module HCB_0 (x, partial_clause, clk, valid);
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= 1'b1;
			partial_clause[0][1] 	= 1'b1;
			partial_clause[0][2] 	= 1'b1;
			partial_clause[0][3] 	= 1'b1;
			partial_clause[0][4] 	= 1'b1;
			partial_clause[0][5] 	= 1'b1;
			partial_clause[0][6] 	= 1'b1;
			partial_clause[0][7] 	= 1'b0;
			partial_clause[0][8] 	= 1'b1;
			partial_clause[0][9] 	= 1'b0;
			partial_clause[0][10] 	= 1'b1;
			partial_clause[0][11] 	= 1'b1;
			partial_clause[0][12] 	= 1'b0;
			partial_clause[0][13] 	= 1'b1;
			partial_clause[0][14] 	= 1'b1;
			partial_clause[0][15] 	= 1'b1;
			partial_clause[0][16] 	= 1'b1;
			partial_clause[0][17] 	= 1'b1;
			partial_clause[0][18] 	= 1'b1;
			partial_clause[0][19] 	= 1'b1;
			partial_clause[0][20] 	= 1'b1;
			partial_clause[0][21] 	= 1'b1;
			partial_clause[0][22] 	= 1'b1;
			partial_clause[0][23] 	= 1'b1;
			partial_clause[0][24] 	= 1'b1;
			partial_clause[0][25] 	= 1'b1;
			partial_clause[0][26] 	= 1'b1;
			partial_clause[0][27] 	= 1'b1;
			partial_clause[0][28] 	= 1'b1;
			partial_clause[0][29] 	= 1'b1;
			partial_clause[0][30] 	= 1'b1;
			partial_clause[0][31] 	= x[54];
			partial_clause[0][32] 	= 1'b1;
			partial_clause[0][33] 	= 1'b0;
			partial_clause[0][34] 	= 1'b1;
			partial_clause[0][35] 	= 1'b1;
			partial_clause[0][36] 	= 1'b1;
			partial_clause[0][37] 	= 1'b1;
			partial_clause[0][38] 	= 1'b1;
			partial_clause[0][39] 	= 1'b1;
			partial_clause[0][40] 	= 1'b1;
			partial_clause[0][41] 	= 1'b1;
			partial_clause[0][42] 	= 1'b0;
			partial_clause[0][43] 	= 1'b1;
			partial_clause[0][44] 	= 1'b1;
			partial_clause[0][45] 	= 1'b1;
			partial_clause[0][46] 	= 1'b1;
			partial_clause[0][47] 	= 1'b1;
			partial_clause[0][48] 	= 1'b1;
			partial_clause[0][49] 	= 1'b1;
			partial_clause[0][50] 	= 1'b1;
			partial_clause[0][51] 	= 1'b1;
			partial_clause[0][52] 	= x[3];
			partial_clause[0][53] 	= 1'b1;
			partial_clause[0][54] 	= 1'b1;
			partial_clause[0][55] 	= 1'b1;
			partial_clause[0][56] 	= 1'b1;
			partial_clause[0][57] 	= 1'b0;
			partial_clause[0][58] 	= 1'b1;
			partial_clause[0][59] 	= x[53];
			partial_clause[0][60] 	= 1'b1;
			partial_clause[0][61] 	= x[34];
			partial_clause[0][62] 	= 1'b1;
			partial_clause[0][63] 	= 1'b1;
			partial_clause[0][64] 	= 1'b1;
			partial_clause[0][65] 	= 1'b1;
			partial_clause[0][66] 	= 1'b0;
			partial_clause[0][67] 	= 1'b1;
			partial_clause[0][68] 	= 1'b0;
			partial_clause[0][69] 	= 1'b1;
			partial_clause[0][70] 	= 1'b1;
			partial_clause[0][71] 	= 1'b1;
			partial_clause[0][72] 	= 1'b1;
			partial_clause[0][73] 	= 1'b1;
			partial_clause[0][74] 	= 1'b1;
			partial_clause[0][75] 	= x[53];
			partial_clause[0][76] 	= x[1];
			partial_clause[0][77] 	= 1'b1;
			partial_clause[0][78] 	= 1'b1;
			partial_clause[0][79] 	= 1'b1;
			partial_clause[0][80] 	= x[0];
			partial_clause[0][81] 	= 1'b1;
			partial_clause[0][82] 	= 1'b1;
			partial_clause[0][83] 	= 1'b1;
			partial_clause[0][84] 	= 1'b1;
			partial_clause[0][85] 	= 1'b1;
			partial_clause[0][86] 	= 1'b1;
			partial_clause[0][87] 	= 1'b0;
			partial_clause[0][88] 	= 1'b1;
			partial_clause[0][89] 	= 1'b1;
			partial_clause[0][90] 	= 1'b1;
			partial_clause[0][91] 	= 1'b1;
			partial_clause[0][92] 	= 1'b1;
			partial_clause[0][93] 	= 1'b1;
			partial_clause[0][94] 	= 1'b1;
			partial_clause[0][95] 	= 1'b1;
			partial_clause[0][96] 	= x[53];
			partial_clause[0][97] 	= 1'b1;
			partial_clause[0][98] 	= 1'b1;
			partial_clause[0][99] 	= 1'b1;
			partial_clause[0][100] 	= 1'b1;
			partial_clause[0][101] 	= 1'b1;
			partial_clause[0][102] 	= ~x[6] & ~x[24];
			partial_clause[0][103] 	= 1'b1;
			partial_clause[0][104] 	= 1'b1;
			partial_clause[0][105] 	= 1'b1;
			partial_clause[0][106] 	= 1'b1;
			partial_clause[0][107] 	= 1'b1;
			partial_clause[0][108] 	= 1'b1;
			partial_clause[0][109] 	= 1'b1;
			partial_clause[0][110] 	= 1'b1;
			partial_clause[0][111] 	= 1'b1;
			partial_clause[0][112] 	= ~x[37] & ~x[38];
			partial_clause[0][113] 	= 1'b1;
			partial_clause[0][114] 	= 1'b1;
			partial_clause[0][115] 	= 1'b1;
			partial_clause[0][116] 	= 1'b1;
			partial_clause[0][117] 	= 1'b1;
			partial_clause[0][118] 	= 1'b1;
			partial_clause[0][119] 	= 1'b1;
			partial_clause[0][120] 	= 1'b1;
			partial_clause[0][121] 	= 1'b1;
			partial_clause[0][122] 	= 1'b0;
			partial_clause[0][123] 	= 1'b1;
			partial_clause[0][124] 	= 1'b1;
			partial_clause[0][125] 	= 1'b1;
			partial_clause[0][126] 	= 1'b1;
			partial_clause[0][127] 	= 1'b1;
			partial_clause[0][128] 	= 1'b1;
			partial_clause[0][129] 	= 1'b1;
			partial_clause[0][130] 	= 1'b1;
			partial_clause[0][131] 	= 1'b1;
			partial_clause[0][132] 	= ~x[5];
			partial_clause[0][133] 	= 1'b1;
			partial_clause[0][134] 	= 1'b1;
			partial_clause[0][135] 	= 1'b1;
			partial_clause[0][136] 	= 1'b1;
			partial_clause[0][137] 	= 1'b0;
			partial_clause[0][138] 	= 1'b1;
			partial_clause[0][139] 	= 1'b1;
			partial_clause[0][140] 	= 1'b1;
			partial_clause[0][141] 	= 1'b1;
			partial_clause[0][142] 	= 1'b1;
			partial_clause[0][143] 	= 1'b1;
			partial_clause[0][144] 	= 1'b1;
			partial_clause[0][145] 	= 1'b1;
			partial_clause[0][146] 	= 1'b1;
			partial_clause[0][147] 	= 1'b1;
			partial_clause[0][148] 	= 1'b1;
			partial_clause[0][149] 	= 1'b1;
			partial_clause[0][150] 	= 1'b1;
			partial_clause[0][151] 	= 1'b1;
			partial_clause[0][152] 	= 1'b1;
			partial_clause[0][153] 	= 1'b1;
			partial_clause[0][154] 	= 1'b0;
			partial_clause[0][155] 	= 1'b1;
			partial_clause[0][156] 	= 1'b1;
			partial_clause[0][157] 	= 1'b1;
			partial_clause[0][158] 	= 1'b1;
			partial_clause[0][159] 	= 1'b1;
			partial_clause[0][160] 	= 1'b1;
			partial_clause[0][161] 	= 1'b1;
			partial_clause[0][162] 	= 1'b1;
			partial_clause[0][163] 	= 1'b1;
			partial_clause[0][164] 	= 1'b1;
			partial_clause[0][165] 	= 1'b1;
			partial_clause[0][166] 	= 1'b1;
			partial_clause[0][167] 	= 1'b1;
			partial_clause[0][168] 	= 1'b1;
			partial_clause[0][169] 	= 1'b1;
			partial_clause[0][170] 	= 1'b1;
			partial_clause[0][171] 	= 1'b1;
			partial_clause[0][172] 	= 1'b1;
			partial_clause[0][173] 	= 1'b1;
			partial_clause[0][174] 	= 1'b1;
			partial_clause[0][175] 	= 1'b1;
			partial_clause[0][176] 	= 1'b1;
			partial_clause[0][177] 	= 1'b1;
			partial_clause[0][178] 	= 1'b1;
			partial_clause[0][179] 	= 1'b1;
			partial_clause[0][180] 	= 1'b1;
			partial_clause[0][181] 	= 1'b1;
			partial_clause[0][182] 	= 1'b1;
			partial_clause[0][183] 	= 1'b1;
			partial_clause[0][184] 	= 1'b1;
			partial_clause[0][185] 	= 1'b1;
			partial_clause[0][186] 	= 1'b1;
			partial_clause[0][187] 	= 1'b1;
			partial_clause[0][188] 	= 1'b1;
			partial_clause[0][189] 	= 1'b1;
			partial_clause[0][190] 	= 1'b1;
			partial_clause[0][191] 	= 1'b1;
			partial_clause[0][192] 	= 1'b1;
			partial_clause[0][193] 	= 1'b1;
			partial_clause[0][194] 	= 1'b1;
			partial_clause[0][195] 	= 1'b1;
			partial_clause[0][196] 	= 1'b1;
			partial_clause[0][197] 	= 1'b1;
			partial_clause[0][198] 	= 1'b1;
			partial_clause[0][199] 	= 1'b1;
			// Class 1
			partial_clause[1][0] 	= 1'b1;
			partial_clause[1][1] 	= 1'b1;
			partial_clause[1][2] 	= 1'b1;
			partial_clause[1][3] 	= 1'b1;
			partial_clause[1][4] 	= 1'b1;
			partial_clause[1][5] 	= 1'b1;
			partial_clause[1][6] 	= x[3];
			partial_clause[1][7] 	= 1'b1;
			partial_clause[1][8] 	= 1'b1;
			partial_clause[1][9] 	= 1'b1;
			partial_clause[1][10] 	= 1'b1;
			partial_clause[1][11] 	= 1'b1;
			partial_clause[1][12] 	= 1'b1;
			partial_clause[1][13] 	= 1'b1;
			partial_clause[1][14] 	= 1'b1;
			partial_clause[1][15] 	= 1'b1;
			partial_clause[1][16] 	= 1'b0;
			partial_clause[1][17] 	= 1'b0;
			partial_clause[1][18] 	= x[2];
			partial_clause[1][19] 	= 1'b1;
			partial_clause[1][20] 	= 1'b0;
			partial_clause[1][21] 	= 1'b1;
			partial_clause[1][22] 	= 1'b1;
			partial_clause[1][23] 	= 1'b0;
			partial_clause[1][24] 	= 1'b1;
			partial_clause[1][25] 	= 1'b1;
			partial_clause[1][26] 	= 1'b1;
			partial_clause[1][27] 	= 1'b1;
			partial_clause[1][28] 	= x[16];
			partial_clause[1][29] 	= 1'b1;
			partial_clause[1][30] 	= 1'b1;
			partial_clause[1][31] 	= 1'b1;
			partial_clause[1][32] 	= x[23];
			partial_clause[1][33] 	= 1'b1;
			partial_clause[1][34] 	= 1'b1;
			partial_clause[1][35] 	= 1'b1;
			partial_clause[1][36] 	= 1'b1;
			partial_clause[1][37] 	= 1'b1;
			partial_clause[1][38] 	= 1'b1;
			partial_clause[1][39] 	= 1'b1;
			partial_clause[1][40] 	= 1'b1;
			partial_clause[1][41] 	= 1'b1;
			partial_clause[1][42] 	= 1'b1;
			partial_clause[1][43] 	= 1'b1;
			partial_clause[1][44] 	= 1'b0;
			partial_clause[1][45] 	= 1'b1;
			partial_clause[1][46] 	= 1'b1;
			partial_clause[1][47] 	= 1'b1;
			partial_clause[1][48] 	= x[6];
			partial_clause[1][49] 	= 1'b1;
			partial_clause[1][50] 	= x[10];
			partial_clause[1][51] 	= 1'b1;
			partial_clause[1][52] 	= 1'b1;
			partial_clause[1][53] 	= x[26];
			partial_clause[1][54] 	= 1'b1;
			partial_clause[1][55] 	= 1'b1;
			partial_clause[1][56] 	= x[46];
			partial_clause[1][57] 	= 1'b1;
			partial_clause[1][58] 	= 1'b1;
			partial_clause[1][59] 	= 1'b1;
			partial_clause[1][60] 	= 1'b1;
			partial_clause[1][61] 	= 1'b0;
			partial_clause[1][62] 	= 1'b1;
			partial_clause[1][63] 	= 1'b1;
			partial_clause[1][64] 	= 1'b1;
			partial_clause[1][65] 	= 1'b1;
			partial_clause[1][66] 	= 1'b1;
			partial_clause[1][67] 	= 1'b1;
			partial_clause[1][68] 	= 1'b1;
			partial_clause[1][69] 	= x[38];
			partial_clause[1][70] 	= 1'b1;
			partial_clause[1][71] 	= 1'b1;
			partial_clause[1][72] 	= 1'b1;
			partial_clause[1][73] 	= 1'b1;
			partial_clause[1][74] 	= 1'b1;
			partial_clause[1][75] 	= 1'b1;
			partial_clause[1][76] 	= 1'b1;
			partial_clause[1][77] 	= 1'b1;
			partial_clause[1][78] 	= 1'b1;
			partial_clause[1][79] 	= 1'b1;
			partial_clause[1][80] 	= 1'b1;
			partial_clause[1][81] 	= 1'b0;
			partial_clause[1][82] 	= x[44];
			partial_clause[1][83] 	= 1'b0;
			partial_clause[1][84] 	= 1'b1;
			partial_clause[1][85] 	= 1'b1;
			partial_clause[1][86] 	= x[39];
			partial_clause[1][87] 	= 1'b1;
			partial_clause[1][88] 	= x[17];
			partial_clause[1][89] 	= 1'b1;
			partial_clause[1][90] 	= 1'b1;
			partial_clause[1][91] 	= 1'b1;
			partial_clause[1][92] 	= 1'b1;
			partial_clause[1][93] 	= 1'b0;
			partial_clause[1][94] 	= 1'b1;
			partial_clause[1][95] 	= 1'b1;
			partial_clause[1][96] 	= 1'b0;
			partial_clause[1][97] 	= 1'b1;
			partial_clause[1][98] 	= 1'b1;
			partial_clause[1][99] 	= 1'b1;
			partial_clause[1][100] 	= 1'b1;
			partial_clause[1][101] 	= 1'b1;
			partial_clause[1][102] 	= 1'b1;
			partial_clause[1][103] 	= 1'b1;
			partial_clause[1][104] 	= 1'b1;
			partial_clause[1][105] 	= 1'b1;
			partial_clause[1][106] 	= 1'b1;
			partial_clause[1][107] 	= 1'b1;
			partial_clause[1][108] 	= 1'b0;
			partial_clause[1][109] 	= 1'b1;
			partial_clause[1][110] 	= 1'b1;
			partial_clause[1][111] 	= 1'b1;
			partial_clause[1][112] 	= 1'b1;
			partial_clause[1][113] 	= 1'b1;
			partial_clause[1][114] 	= 1'b1;
			partial_clause[1][115] 	= 1'b1;
			partial_clause[1][116] 	= 1'b1;
			partial_clause[1][117] 	= 1'b0;
			partial_clause[1][118] 	= 1'b1;
			partial_clause[1][119] 	= 1'b1;
			partial_clause[1][120] 	= 1'b1;
			partial_clause[1][121] 	= 1'b1;
			partial_clause[1][122] 	= 1'b1;
			partial_clause[1][123] 	= 1'b1;
			partial_clause[1][124] 	= 1'b1;
			partial_clause[1][125] 	= 1'b1;
			partial_clause[1][126] 	= 1'b1;
			partial_clause[1][127] 	= 1'b1;
			partial_clause[1][128] 	= 1'b1;
			partial_clause[1][129] 	= 1'b0;
			partial_clause[1][130] 	= 1'b1;
			partial_clause[1][131] 	= 1'b1;
			partial_clause[1][132] 	= 1'b1;
			partial_clause[1][133] 	= 1'b1;
			partial_clause[1][134] 	= 1'b1;
			partial_clause[1][135] 	= 1'b0;
			partial_clause[1][136] 	= 1'b1;
			partial_clause[1][137] 	= 1'b0;
			partial_clause[1][138] 	= 1'b1;
			partial_clause[1][139] 	= 1'b1;
			partial_clause[1][140] 	= 1'b1;
			partial_clause[1][141] 	= 1'b1;
			partial_clause[1][142] 	= 1'b1;
			partial_clause[1][143] 	= 1'b1;
			partial_clause[1][144] 	= 1'b1;
			partial_clause[1][145] 	= 1'b1;
			partial_clause[1][146] 	= 1'b1;
			partial_clause[1][147] 	= 1'b1;
			partial_clause[1][148] 	= 1'b1;
			partial_clause[1][149] 	= 1'b1;
			partial_clause[1][150] 	= 1'b1;
			partial_clause[1][151] 	= 1'b1;
			partial_clause[1][152] 	= 1'b1;
			partial_clause[1][153] 	= 1'b1;
			partial_clause[1][154] 	= 1'b1;
			partial_clause[1][155] 	= 1'b1;
			partial_clause[1][156] 	= 1'b1;
			partial_clause[1][157] 	= 1'b1;
			partial_clause[1][158] 	= 1'b1;
			partial_clause[1][159] 	= 1'b1;
			partial_clause[1][160] 	= 1'b1;
			partial_clause[1][161] 	= 1'b1;
			partial_clause[1][162] 	= 1'b1;
			partial_clause[1][163] 	= 1'b1;
			partial_clause[1][164] 	= 1'b0;
			partial_clause[1][165] 	= 1'b1;
			partial_clause[1][166] 	= 1'b1;
			partial_clause[1][167] 	= 1'b1;
			partial_clause[1][168] 	= 1'b1;
			partial_clause[1][169] 	= 1'b1;
			partial_clause[1][170] 	= 1'b1;
			partial_clause[1][171] 	= 1'b1;
			partial_clause[1][172] 	= 1'b1;
			partial_clause[1][173] 	= 1'b1;
			partial_clause[1][174] 	= 1'b1;
			partial_clause[1][175] 	= 1'b1;
			partial_clause[1][176] 	= 1'b1;
			partial_clause[1][177] 	= 1'b1;
			partial_clause[1][178] 	= 1'b1;
			partial_clause[1][179] 	= 1'b1;
			partial_clause[1][180] 	= 1'b1;
			partial_clause[1][181] 	= 1'b1;
			partial_clause[1][182] 	= 1'b1;
			partial_clause[1][183] 	= 1'b1;
			partial_clause[1][184] 	= 1'b1;
			partial_clause[1][185] 	= 1'b0;
			partial_clause[1][186] 	= 1'b1;
			partial_clause[1][187] 	= 1'b1;
			partial_clause[1][188] 	= 1'b1;
			partial_clause[1][189] 	= 1'b1;
			partial_clause[1][190] 	= 1'b0;
			partial_clause[1][191] 	= 1'b1;
			partial_clause[1][192] 	= 1'b1;
			partial_clause[1][193] 	= 1'b1;
			partial_clause[1][194] 	= 1'b1;
			partial_clause[1][195] 	= 1'b1;
			partial_clause[1][196] 	= 1'b1;
			partial_clause[1][197] 	= 1'b1;
			partial_clause[1][198] 	= 1'b1;
			partial_clause[1][199] 	= 1'b1;
			// Class 2
			partial_clause[2][0] 	= 1'b1;
			partial_clause[2][1] 	= 1'b1;
			partial_clause[2][2] 	= 1'b1;
			partial_clause[2][3] 	= 1'b1;
			partial_clause[2][4] 	= 1'b1;
			partial_clause[2][5] 	= x[8];
			partial_clause[2][6] 	= 1'b1;
			partial_clause[2][7] 	= 1'b1;
			partial_clause[2][8] 	= 1'b1;
			partial_clause[2][9] 	= 1'b1;
			partial_clause[2][10] 	= 1'b1;
			partial_clause[2][11] 	= 1'b1;
			partial_clause[2][12] 	= 1'b1;
			partial_clause[2][13] 	= 1'b1;
			partial_clause[2][14] 	= 1'b1;
			partial_clause[2][15] 	= x[41];
			partial_clause[2][16] 	= 1'b1;
			partial_clause[2][17] 	= 1'b1;
			partial_clause[2][18] 	= 1'b1;
			partial_clause[2][19] 	= 1'b1;
			partial_clause[2][20] 	= 1'b1;
			partial_clause[2][21] 	= 1'b1;
			partial_clause[2][22] 	= 1'b1;
			partial_clause[2][23] 	= 1'b1;
			partial_clause[2][24] 	= 1'b1;
			partial_clause[2][25] 	= 1'b1;
			partial_clause[2][26] 	= 1'b1;
			partial_clause[2][27] 	= 1'b1;
			partial_clause[2][28] 	= 1'b1;
			partial_clause[2][29] 	= 1'b1;
			partial_clause[2][30] 	= 1'b0;
			partial_clause[2][31] 	= 1'b1;
			partial_clause[2][32] 	= 1'b1;
			partial_clause[2][33] 	= 1'b1;
			partial_clause[2][34] 	= 1'b1;
			partial_clause[2][35] 	= 1'b1;
			partial_clause[2][36] 	= 1'b1;
			partial_clause[2][37] 	= 1'b1;
			partial_clause[2][38] 	= 1'b1;
			partial_clause[2][39] 	= 1'b1;
			partial_clause[2][40] 	= 1'b1;
			partial_clause[2][41] 	= 1'b1;
			partial_clause[2][42] 	= 1'b1;
			partial_clause[2][43] 	= 1'b1;
			partial_clause[2][44] 	= 1'b1;
			partial_clause[2][45] 	= 1'b1;
			partial_clause[2][46] 	= 1'b1;
			partial_clause[2][47] 	= 1'b1;
			partial_clause[2][48] 	= 1'b1;
			partial_clause[2][49] 	= x[11];
			partial_clause[2][50] 	= 1'b1;
			partial_clause[2][51] 	= 1'b1;
			partial_clause[2][52] 	= 1'b1;
			partial_clause[2][53] 	= 1'b1;
			partial_clause[2][54] 	= 1'b1;
			partial_clause[2][55] 	= 1'b1;
			partial_clause[2][56] 	= 1'b1;
			partial_clause[2][57] 	= 1'b1;
			partial_clause[2][58] 	= 1'b1;
			partial_clause[2][59] 	= 1'b1;
			partial_clause[2][60] 	= 1'b1;
			partial_clause[2][61] 	= 1'b1;
			partial_clause[2][62] 	= 1'b1;
			partial_clause[2][63] 	= 1'b1;
			partial_clause[2][64] 	= 1'b1;
			partial_clause[2][65] 	= 1'b1;
			partial_clause[2][66] 	= 1'b1;
			partial_clause[2][67] 	= 1'b1;
			partial_clause[2][68] 	= 1'b1;
			partial_clause[2][69] 	= 1'b1;
			partial_clause[2][70] 	= 1'b1;
			partial_clause[2][71] 	= 1'b1;
			partial_clause[2][72] 	= 1'b1;
			partial_clause[2][73] 	= 1'b0;
			partial_clause[2][74] 	= 1'b1;
			partial_clause[2][75] 	= 1'b1;
			partial_clause[2][76] 	= 1'b1;
			partial_clause[2][77] 	= 1'b1;
			partial_clause[2][78] 	= 1'b1;
			partial_clause[2][79] 	= 1'b1;
			partial_clause[2][80] 	= 1'b1;
			partial_clause[2][81] 	= 1'b1;
			partial_clause[2][82] 	= 1'b1;
			partial_clause[2][83] 	= 1'b1;
			partial_clause[2][84] 	= 1'b1;
			partial_clause[2][85] 	= 1'b1;
			partial_clause[2][86] 	= 1'b1;
			partial_clause[2][87] 	= 1'b1;
			partial_clause[2][88] 	= x[14];
			partial_clause[2][89] 	= 1'b1;
			partial_clause[2][90] 	= 1'b1;
			partial_clause[2][91] 	= 1'b1;
			partial_clause[2][92] 	= 1'b1;
			partial_clause[2][93] 	= 1'b1;
			partial_clause[2][94] 	= 1'b1;
			partial_clause[2][95] 	= 1'b1;
			partial_clause[2][96] 	= 1'b1;
			partial_clause[2][97] 	= 1'b1;
			partial_clause[2][98] 	= 1'b1;
			partial_clause[2][99] 	= 1'b1;
			partial_clause[2][100] 	= 1'b1;
			partial_clause[2][101] 	= 1'b0;
			partial_clause[2][102] 	= ~x[60];
			partial_clause[2][103] 	= 1'b1;
			partial_clause[2][104] 	= 1'b1;
			partial_clause[2][105] 	= 1'b1;
			partial_clause[2][106] 	= 1'b0;
			partial_clause[2][107] 	= 1'b1;
			partial_clause[2][108] 	= 1'b1;
			partial_clause[2][109] 	= 1'b1;
			partial_clause[2][110] 	= 1'b1;
			partial_clause[2][111] 	= 1'b1;
			partial_clause[2][112] 	= 1'b1;
			partial_clause[2][113] 	= 1'b0;
			partial_clause[2][114] 	= 1'b1;
			partial_clause[2][115] 	= 1'b1;
			partial_clause[2][116] 	= 1'b0;
			partial_clause[2][117] 	= 1'b1;
			partial_clause[2][118] 	= 1'b1;
			partial_clause[2][119] 	= 1'b1;
			partial_clause[2][120] 	= 1'b1;
			partial_clause[2][121] 	= 1'b1;
			partial_clause[2][122] 	= 1'b1;
			partial_clause[2][123] 	= 1'b1;
			partial_clause[2][124] 	= 1'b0;
			partial_clause[2][125] 	= 1'b1;
			partial_clause[2][126] 	= 1'b1;
			partial_clause[2][127] 	= 1'b1;
			partial_clause[2][128] 	= 1'b1;
			partial_clause[2][129] 	= 1'b1;
			partial_clause[2][130] 	= 1'b1;
			partial_clause[2][131] 	= 1'b1;
			partial_clause[2][132] 	= 1'b1;
			partial_clause[2][133] 	= 1'b1;
			partial_clause[2][134] 	= 1'b1;
			partial_clause[2][135] 	= 1'b0;
			partial_clause[2][136] 	= 1'b1;
			partial_clause[2][137] 	= 1'b1;
			partial_clause[2][138] 	= 1'b1;
			partial_clause[2][139] 	= 1'b1;
			partial_clause[2][140] 	= 1'b1;
			partial_clause[2][141] 	= 1'b1;
			partial_clause[2][142] 	= 1'b1;
			partial_clause[2][143] 	= 1'b1;
			partial_clause[2][144] 	= 1'b1;
			partial_clause[2][145] 	= 1'b1;
			partial_clause[2][146] 	= 1'b1;
			partial_clause[2][147] 	= 1'b1;
			partial_clause[2][148] 	= ~x[48];
			partial_clause[2][149] 	= 1'b1;
			partial_clause[2][150] 	= 1'b1;
			partial_clause[2][151] 	= 1'b1;
			partial_clause[2][152] 	= 1'b1;
			partial_clause[2][153] 	= 1'b1;
			partial_clause[2][154] 	= 1'b0;
			partial_clause[2][155] 	= 1'b1;
			partial_clause[2][156] 	= 1'b1;
			partial_clause[2][157] 	= 1'b1;
			partial_clause[2][158] 	= 1'b1;
			partial_clause[2][159] 	= 1'b1;
			partial_clause[2][160] 	= 1'b1;
			partial_clause[2][161] 	= 1'b1;
			partial_clause[2][162] 	= 1'b1;
			partial_clause[2][163] 	= 1'b1;
			partial_clause[2][164] 	= 1'b1;
			partial_clause[2][165] 	= 1'b1;
			partial_clause[2][166] 	= 1'b1;
			partial_clause[2][167] 	= 1'b1;
			partial_clause[2][168] 	= 1'b1;
			partial_clause[2][169] 	= 1'b1;
			partial_clause[2][170] 	= 1'b0;
			partial_clause[2][171] 	= x[56];
			partial_clause[2][172] 	= 1'b1;
			partial_clause[2][173] 	= 1'b1;
			partial_clause[2][174] 	= 1'b1;
			partial_clause[2][175] 	= 1'b1;
			partial_clause[2][176] 	= 1'b1;
			partial_clause[2][177] 	= 1'b1;
			partial_clause[2][178] 	= 1'b1;
			partial_clause[2][179] 	= 1'b0;
			partial_clause[2][180] 	= 1'b1;
			partial_clause[2][181] 	= 1'b1;
			partial_clause[2][182] 	= 1'b1;
			partial_clause[2][183] 	= 1'b1;
			partial_clause[2][184] 	= 1'b0;
			partial_clause[2][185] 	= 1'b1;
			partial_clause[2][186] 	= 1'b1;
			partial_clause[2][187] 	= 1'b1;
			partial_clause[2][188] 	= 1'b0;
			partial_clause[2][189] 	= 1'b1;
			partial_clause[2][190] 	= 1'b1;
			partial_clause[2][191] 	= 1'b1;
			partial_clause[2][192] 	= 1'b1;
			partial_clause[2][193] 	= 1'b1;
			partial_clause[2][194] 	= 1'b1;
			partial_clause[2][195] 	= 1'b1;
			partial_clause[2][196] 	= 1'b1;
			partial_clause[2][197] 	= 1'b1;
			partial_clause[2][198] 	= 1'b1;
			partial_clause[2][199] 	= 1'b1;
			// Class 3
			partial_clause[3][0] 	= 1'b1;
			partial_clause[3][1] 	= 1'b1;
			partial_clause[3][2] 	= 1'b1;
			partial_clause[3][3] 	= 1'b1;
			partial_clause[3][4] 	= 1'b1;
			partial_clause[3][5] 	= 1'b1;
			partial_clause[3][6] 	= 1'b0;
			partial_clause[3][7] 	= 1'b1;
			partial_clause[3][8] 	= 1'b1;
			partial_clause[3][9] 	= 1'b1;
			partial_clause[3][10] 	= 1'b1;
			partial_clause[3][11] 	= 1'b1;
			partial_clause[3][12] 	= 1'b0;
			partial_clause[3][13] 	= 1'b1;
			partial_clause[3][14] 	= x[36];
			partial_clause[3][15] 	= 1'b1;
			partial_clause[3][16] 	= 1'b1;
			partial_clause[3][17] 	= 1'b1;
			partial_clause[3][18] 	= 1'b1;
			partial_clause[3][19] 	= 1'b1;
			partial_clause[3][20] 	= 1'b1;
			partial_clause[3][21] 	= 1'b1;
			partial_clause[3][22] 	= 1'b0;
			partial_clause[3][23] 	= 1'b1;
			partial_clause[3][24] 	= 1'b1;
			partial_clause[3][25] 	= 1'b1;
			partial_clause[3][26] 	= x[1];
			partial_clause[3][27] 	= 1'b1;
			partial_clause[3][28] 	= 1'b1;
			partial_clause[3][29] 	= 1'b1;
			partial_clause[3][30] 	= 1'b1;
			partial_clause[3][31] 	= 1'b1;
			partial_clause[3][32] 	= 1'b1;
			partial_clause[3][33] 	= 1'b1;
			partial_clause[3][34] 	= 1'b1;
			partial_clause[3][35] 	= 1'b1;
			partial_clause[3][36] 	= 1'b1;
			partial_clause[3][37] 	= 1'b1;
			partial_clause[3][38] 	= 1'b1;
			partial_clause[3][39] 	= 1'b1;
			partial_clause[3][40] 	= 1'b1;
			partial_clause[3][41] 	= ~x[40];
			partial_clause[3][42] 	= 1'b1;
			partial_clause[3][43] 	= 1'b1;
			partial_clause[3][44] 	= 1'b1;
			partial_clause[3][45] 	= 1'b0;
			partial_clause[3][46] 	= 1'b1;
			partial_clause[3][47] 	= 1'b1;
			partial_clause[3][48] 	= 1'b1;
			partial_clause[3][49] 	= 1'b1;
			partial_clause[3][50] 	= 1'b1;
			partial_clause[3][51] 	= 1'b1;
			partial_clause[3][52] 	= 1'b1;
			partial_clause[3][53] 	= 1'b1;
			partial_clause[3][54] 	= 1'b1;
			partial_clause[3][55] 	= 1'b1;
			partial_clause[3][56] 	= 1'b1;
			partial_clause[3][57] 	= 1'b1;
			partial_clause[3][58] 	= 1'b1;
			partial_clause[3][59] 	= 1'b1;
			partial_clause[3][60] 	= 1'b1;
			partial_clause[3][61] 	= 1'b1;
			partial_clause[3][62] 	= 1'b1;
			partial_clause[3][63] 	= 1'b1;
			partial_clause[3][64] 	= 1'b1;
			partial_clause[3][65] 	= 1'b1;
			partial_clause[3][66] 	= 1'b1;
			partial_clause[3][67] 	= 1'b0;
			partial_clause[3][68] 	= 1'b1;
			partial_clause[3][69] 	= 1'b1;
			partial_clause[3][70] 	= 1'b1;
			partial_clause[3][71] 	= 1'b1;
			partial_clause[3][72] 	= 1'b0;
			partial_clause[3][73] 	= x[0];
			partial_clause[3][74] 	= 1'b1;
			partial_clause[3][75] 	= 1'b1;
			partial_clause[3][76] 	= 1'b1;
			partial_clause[3][77] 	= 1'b1;
			partial_clause[3][78] 	= 1'b1;
			partial_clause[3][79] 	= 1'b1;
			partial_clause[3][80] 	= 1'b1;
			partial_clause[3][81] 	= 1'b1;
			partial_clause[3][82] 	= x[34];
			partial_clause[3][83] 	= 1'b1;
			partial_clause[3][84] 	= 1'b0;
			partial_clause[3][85] 	= x[30];
			partial_clause[3][86] 	= 1'b1;
			partial_clause[3][87] 	= 1'b1;
			partial_clause[3][88] 	= 1'b1;
			partial_clause[3][89] 	= 1'b1;
			partial_clause[3][90] 	= 1'b1;
			partial_clause[3][91] 	= 1'b0;
			partial_clause[3][92] 	= 1'b1;
			partial_clause[3][93] 	= 1'b1;
			partial_clause[3][94] 	= 1'b1;
			partial_clause[3][95] 	= 1'b1;
			partial_clause[3][96] 	= 1'b1;
			partial_clause[3][97] 	= 1'b1;
			partial_clause[3][98] 	= 1'b1;
			partial_clause[3][99] 	= 1'b1;
			partial_clause[3][100] 	= 1'b1;
			partial_clause[3][101] 	= 1'b1;
			partial_clause[3][102] 	= 1'b1;
			partial_clause[3][103] 	= 1'b1;
			partial_clause[3][104] 	= 1'b1;
			partial_clause[3][105] 	= 1'b1;
			partial_clause[3][106] 	= 1'b1;
			partial_clause[3][107] 	= 1'b1;
			partial_clause[3][108] 	= 1'b1;
			partial_clause[3][109] 	= 1'b1;
			partial_clause[3][110] 	= 1'b1;
			partial_clause[3][111] 	= 1'b0;
			partial_clause[3][112] 	= 1'b1;
			partial_clause[3][113] 	= 1'b1;
			partial_clause[3][114] 	= 1'b1;
			partial_clause[3][115] 	= 1'b1;
			partial_clause[3][116] 	= 1'b1;
			partial_clause[3][117] 	= 1'b1;
			partial_clause[3][118] 	= 1'b1;
			partial_clause[3][119] 	= 1'b1;
			partial_clause[3][120] 	= 1'b1;
			partial_clause[3][121] 	= 1'b1;
			partial_clause[3][122] 	= 1'b1;
			partial_clause[3][123] 	= 1'b1;
			partial_clause[3][124] 	= 1'b1;
			partial_clause[3][125] 	= 1'b1;
			partial_clause[3][126] 	= 1'b1;
			partial_clause[3][127] 	= 1'b1;
			partial_clause[3][128] 	= 1'b1;
			partial_clause[3][129] 	= 1'b1;
			partial_clause[3][130] 	= x[25];
			partial_clause[3][131] 	= 1'b1;
			partial_clause[3][132] 	= 1'b1;
			partial_clause[3][133] 	= 1'b1;
			partial_clause[3][134] 	= 1'b1;
			partial_clause[3][135] 	= 1'b1;
			partial_clause[3][136] 	= 1'b1;
			partial_clause[3][137] 	= 1'b1;
			partial_clause[3][138] 	= 1'b1;
			partial_clause[3][139] 	= 1'b1;
			partial_clause[3][140] 	= 1'b1;
			partial_clause[3][141] 	= 1'b1;
			partial_clause[3][142] 	= 1'b1;
			partial_clause[3][143] 	= 1'b0;
			partial_clause[3][144] 	= 1'b1;
			partial_clause[3][145] 	= 1'b1;
			partial_clause[3][146] 	= 1'b1;
			partial_clause[3][147] 	= 1'b1;
			partial_clause[3][148] 	= 1'b1;
			partial_clause[3][149] 	= 1'b1;
			partial_clause[3][150] 	= 1'b1;
			partial_clause[3][151] 	= 1'b1;
			partial_clause[3][152] 	= 1'b1;
			partial_clause[3][153] 	= 1'b1;
			partial_clause[3][154] 	= 1'b1;
			partial_clause[3][155] 	= 1'b1;
			partial_clause[3][156] 	= 1'b1;
			partial_clause[3][157] 	= 1'b1;
			partial_clause[3][158] 	= 1'b1;
			partial_clause[3][159] 	= 1'b1;
			partial_clause[3][160] 	= 1'b1;
			partial_clause[3][161] 	= 1'b1;
			partial_clause[3][162] 	= 1'b1;
			partial_clause[3][163] 	= 1'b1;
			partial_clause[3][164] 	= 1'b1;
			partial_clause[3][165] 	= 1'b1;
			partial_clause[3][166] 	= 1'b1;
			partial_clause[3][167] 	= 1'b1;
			partial_clause[3][168] 	= 1'b0;
			partial_clause[3][169] 	= 1'b1;
			partial_clause[3][170] 	= 1'b1;
			partial_clause[3][171] 	= 1'b1;
			partial_clause[3][172] 	= 1'b1;
			partial_clause[3][173] 	= 1'b1;
			partial_clause[3][174] 	= 1'b1;
			partial_clause[3][175] 	= 1'b1;
			partial_clause[3][176] 	= 1'b1;
			partial_clause[3][177] 	= 1'b1;
			partial_clause[3][178] 	= 1'b0;
			partial_clause[3][179] 	= 1'b1;
			partial_clause[3][180] 	= 1'b1;
			partial_clause[3][181] 	= 1'b0;
			partial_clause[3][182] 	= 1'b1;
			partial_clause[3][183] 	= 1'b1;
			partial_clause[3][184] 	= 1'b1;
			partial_clause[3][185] 	= 1'b1;
			partial_clause[3][186] 	= 1'b1;
			partial_clause[3][187] 	= 1'b1;
			partial_clause[3][188] 	= 1'b1;
			partial_clause[3][189] 	= 1'b1;
			partial_clause[3][190] 	= 1'b1;
			partial_clause[3][191] 	= 1'b1;
			partial_clause[3][192] 	= 1'b1;
			partial_clause[3][193] 	= 1'b1;
			partial_clause[3][194] 	= 1'b1;
			partial_clause[3][195] 	= 1'b1;
			partial_clause[3][196] 	= 1'b1;
			partial_clause[3][197] 	= 1'b1;
			partial_clause[3][198] 	= 1'b1;
			partial_clause[3][199] 	= 1'b1;
			// Class 4
			partial_clause[4][0] 	= 1'b1;
			partial_clause[4][1] 	= 1'b1;
			partial_clause[4][2] 	= 1'b1;
			partial_clause[4][3] 	= 1'b1;
			partial_clause[4][4] 	= 1'b0;
			partial_clause[4][5] 	= 1'b1;
			partial_clause[4][6] 	= 1'b1;
			partial_clause[4][7] 	= x[14];
			partial_clause[4][8] 	= 1'b1;
			partial_clause[4][9] 	= 1'b1;
			partial_clause[4][10] 	= 1'b1;
			partial_clause[4][11] 	= 1'b1;
			partial_clause[4][12] 	= 1'b1;
			partial_clause[4][13] 	= 1'b1;
			partial_clause[4][14] 	= 1'b0;
			partial_clause[4][15] 	= 1'b1;
			partial_clause[4][16] 	= 1'b1;
			partial_clause[4][17] 	= 1'b0;
			partial_clause[4][18] 	= 1'b0;
			partial_clause[4][19] 	= 1'b1;
			partial_clause[4][20] 	= 1'b1;
			partial_clause[4][21] 	= 1'b1;
			partial_clause[4][22] 	= 1'b1;
			partial_clause[4][23] 	= 1'b1;
			partial_clause[4][24] 	= 1'b1;
			partial_clause[4][25] 	= 1'b1;
			partial_clause[4][26] 	= 1'b1;
			partial_clause[4][27] 	= 1'b0;
			partial_clause[4][28] 	= 1'b1;
			partial_clause[4][29] 	= x[9];
			partial_clause[4][30] 	= 1'b1;
			partial_clause[4][31] 	= 1'b1;
			partial_clause[4][32] 	= 1'b1;
			partial_clause[4][33] 	= 1'b0;
			partial_clause[4][34] 	= 1'b1;
			partial_clause[4][35] 	= 1'b1;
			partial_clause[4][36] 	= 1'b1;
			partial_clause[4][37] 	= 1'b0;
			partial_clause[4][38] 	= 1'b1;
			partial_clause[4][39] 	= 1'b1;
			partial_clause[4][40] 	= 1'b1;
			partial_clause[4][41] 	= 1'b1;
			partial_clause[4][42] 	= x[51];
			partial_clause[4][43] 	= 1'b0;
			partial_clause[4][44] 	= 1'b1;
			partial_clause[4][45] 	= 1'b0;
			partial_clause[4][46] 	= 1'b1;
			partial_clause[4][47] 	= x[47];
			partial_clause[4][48] 	= 1'b1;
			partial_clause[4][49] 	= 1'b1;
			partial_clause[4][50] 	= 1'b1;
			partial_clause[4][51] 	= 1'b1;
			partial_clause[4][52] 	= 1'b1;
			partial_clause[4][53] 	= 1'b1;
			partial_clause[4][54] 	= 1'b1;
			partial_clause[4][55] 	= 1'b1;
			partial_clause[4][56] 	= 1'b1;
			partial_clause[4][57] 	= 1'b0;
			partial_clause[4][58] 	= 1'b1;
			partial_clause[4][59] 	= 1'b1;
			partial_clause[4][60] 	= 1'b1;
			partial_clause[4][61] 	= 1'b1;
			partial_clause[4][62] 	= 1'b0;
			partial_clause[4][63] 	= 1'b1;
			partial_clause[4][64] 	= 1'b1;
			partial_clause[4][65] 	= 1'b1;
			partial_clause[4][66] 	= 1'b0;
			partial_clause[4][67] 	= 1'b1;
			partial_clause[4][68] 	= 1'b1;
			partial_clause[4][69] 	= 1'b1;
			partial_clause[4][70] 	= x[33];
			partial_clause[4][71] 	= 1'b1;
			partial_clause[4][72] 	= 1'b0;
			partial_clause[4][73] 	= 1'b1;
			partial_clause[4][74] 	= 1'b1;
			partial_clause[4][75] 	= 1'b1;
			partial_clause[4][76] 	= x[9];
			partial_clause[4][77] 	= 1'b1;
			partial_clause[4][78] 	= 1'b1;
			partial_clause[4][79] 	= 1'b1;
			partial_clause[4][80] 	= 1'b1;
			partial_clause[4][81] 	= 1'b1;
			partial_clause[4][82] 	= 1'b1;
			partial_clause[4][83] 	= 1'b1;
			partial_clause[4][84] 	= 1'b1;
			partial_clause[4][85] 	= 1'b1;
			partial_clause[4][86] 	= 1'b1;
			partial_clause[4][87] 	= x[61];
			partial_clause[4][88] 	= 1'b1;
			partial_clause[4][89] 	= x[8];
			partial_clause[4][90] 	= 1'b1;
			partial_clause[4][91] 	= 1'b1;
			partial_clause[4][92] 	= 1'b1;
			partial_clause[4][93] 	= 1'b1;
			partial_clause[4][94] 	= 1'b0;
			partial_clause[4][95] 	= 1'b1;
			partial_clause[4][96] 	= 1'b1;
			partial_clause[4][97] 	= 1'b1;
			partial_clause[4][98] 	= 1'b0;
			partial_clause[4][99] 	= 1'b1;
			partial_clause[4][100] 	= 1'b1;
			partial_clause[4][101] 	= 1'b1;
			partial_clause[4][102] 	= 1'b1;
			partial_clause[4][103] 	= ~x[53];
			partial_clause[4][104] 	= 1'b1;
			partial_clause[4][105] 	= 1'b1;
			partial_clause[4][106] 	= 1'b1;
			partial_clause[4][107] 	= 1'b1;
			partial_clause[4][108] 	= 1'b1;
			partial_clause[4][109] 	= 1'b1;
			partial_clause[4][110] 	= 1'b1;
			partial_clause[4][111] 	= 1'b1;
			partial_clause[4][112] 	= 1'b1;
			partial_clause[4][113] 	= 1'b1;
			partial_clause[4][114] 	= 1'b1;
			partial_clause[4][115] 	= 1'b1;
			partial_clause[4][116] 	= 1'b1;
			partial_clause[4][117] 	= 1'b1;
			partial_clause[4][118] 	= 1'b1;
			partial_clause[4][119] 	= 1'b1;
			partial_clause[4][120] 	= 1'b1;
			partial_clause[4][121] 	= 1'b1;
			partial_clause[4][122] 	= 1'b1;
			partial_clause[4][123] 	= 1'b1;
			partial_clause[4][124] 	= 1'b1;
			partial_clause[4][125] 	= 1'b1;
			partial_clause[4][126] 	= 1'b1;
			partial_clause[4][127] 	= 1'b1;
			partial_clause[4][128] 	= 1'b1;
			partial_clause[4][129] 	= 1'b1;
			partial_clause[4][130] 	= 1'b1;
			partial_clause[4][131] 	= 1'b1;
			partial_clause[4][132] 	= 1'b1;
			partial_clause[4][133] 	= 1'b1;
			partial_clause[4][134] 	= 1'b1;
			partial_clause[4][135] 	= 1'b1;
			partial_clause[4][136] 	= 1'b1;
			partial_clause[4][137] 	= 1'b1;
			partial_clause[4][138] 	= 1'b1;
			partial_clause[4][139] 	= 1'b1;
			partial_clause[4][140] 	= 1'b1;
			partial_clause[4][141] 	= 1'b1;
			partial_clause[4][142] 	= 1'b1;
			partial_clause[4][143] 	= 1'b1;
			partial_clause[4][144] 	= 1'b1;
			partial_clause[4][145] 	= 1'b1;
			partial_clause[4][146] 	= 1'b1;
			partial_clause[4][147] 	= 1'b1;
			partial_clause[4][148] 	= 1'b1;
			partial_clause[4][149] 	= 1'b1;
			partial_clause[4][150] 	= 1'b1;
			partial_clause[4][151] 	= 1'b1;
			partial_clause[4][152] 	= 1'b1;
			partial_clause[4][153] 	= 1'b1;
			partial_clause[4][154] 	= 1'b1;
			partial_clause[4][155] 	= ~x[24];
			partial_clause[4][156] 	= 1'b1;
			partial_clause[4][157] 	= 1'b1;
			partial_clause[4][158] 	= 1'b1;
			partial_clause[4][159] 	= 1'b1;
			partial_clause[4][160] 	= 1'b1;
			partial_clause[4][161] 	= 1'b1;
			partial_clause[4][162] 	= 1'b1;
			partial_clause[4][163] 	= 1'b1;
			partial_clause[4][164] 	= 1'b1;
			partial_clause[4][165] 	= 1'b1;
			partial_clause[4][166] 	= 1'b1;
			partial_clause[4][167] 	= 1'b1;
			partial_clause[4][168] 	= 1'b1;
			partial_clause[4][169] 	= 1'b1;
			partial_clause[4][170] 	= 1'b1;
			partial_clause[4][171] 	= 1'b1;
			partial_clause[4][172] 	= 1'b1;
			partial_clause[4][173] 	= 1'b1;
			partial_clause[4][174] 	= 1'b1;
			partial_clause[4][175] 	= 1'b1;
			partial_clause[4][176] 	= 1'b1;
			partial_clause[4][177] 	= 1'b1;
			partial_clause[4][178] 	= 1'b1;
			partial_clause[4][179] 	= 1'b1;
			partial_clause[4][180] 	= 1'b1;
			partial_clause[4][181] 	= 1'b1;
			partial_clause[4][182] 	= 1'b1;
			partial_clause[4][183] 	= 1'b1;
			partial_clause[4][184] 	= 1'b1;
			partial_clause[4][185] 	= 1'b1;
			partial_clause[4][186] 	= 1'b1;
			partial_clause[4][187] 	= 1'b1;
			partial_clause[4][188] 	= 1'b1;
			partial_clause[4][189] 	= 1'b1;
			partial_clause[4][190] 	= 1'b1;
			partial_clause[4][191] 	= 1'b1;
			partial_clause[4][192] 	= 1'b1;
			partial_clause[4][193] 	= 1'b1;
			partial_clause[4][194] 	= 1'b1;
			partial_clause[4][195] 	= 1'b1;
			partial_clause[4][196] 	= 1'b1;
			partial_clause[4][197] 	= 1'b1;
			partial_clause[4][198] 	= 1'b1;
			partial_clause[4][199] 	= 1'b1;
			// Class 5
			partial_clause[5][0] 	= 1'b1;
			partial_clause[5][1] 	= 1'b0;
			partial_clause[5][2] 	= 1'b1;
			partial_clause[5][3] 	= 1'b1;
			partial_clause[5][4] 	= 1'b1;
			partial_clause[5][5] 	= 1'b1;
			partial_clause[5][6] 	= 1'b1;
			partial_clause[5][7] 	= x[63];
			partial_clause[5][8] 	= 1'b1;
			partial_clause[5][9] 	= 1'b1;
			partial_clause[5][10] 	= 1'b0;
			partial_clause[5][11] 	= 1'b1;
			partial_clause[5][12] 	= 1'b1;
			partial_clause[5][13] 	= 1'b1;
			partial_clause[5][14] 	= 1'b1;
			partial_clause[5][15] 	= 1'b1;
			partial_clause[5][16] 	= 1'b1;
			partial_clause[5][17] 	= 1'b1;
			partial_clause[5][18] 	= 1'b1;
			partial_clause[5][19] 	= 1'b1;
			partial_clause[5][20] 	= 1'b1;
			partial_clause[5][21] 	= 1'b1;
			partial_clause[5][22] 	= 1'b1;
			partial_clause[5][23] 	= 1'b1;
			partial_clause[5][24] 	= 1'b1;
			partial_clause[5][25] 	= 1'b1;
			partial_clause[5][26] 	= 1'b1;
			partial_clause[5][27] 	= 1'b1;
			partial_clause[5][28] 	= 1'b1;
			partial_clause[5][29] 	= 1'b1;
			partial_clause[5][30] 	= 1'b1;
			partial_clause[5][31] 	= 1'b1;
			partial_clause[5][32] 	= 1'b1;
			partial_clause[5][33] 	= x[14];
			partial_clause[5][34] 	= 1'b1;
			partial_clause[5][35] 	= 1'b1;
			partial_clause[5][36] 	= 1'b1;
			partial_clause[5][37] 	= 1'b1;
			partial_clause[5][38] 	= 1'b1;
			partial_clause[5][39] 	= 1'b1;
			partial_clause[5][40] 	= 1'b1;
			partial_clause[5][41] 	= 1'b1;
			partial_clause[5][42] 	= 1'b1;
			partial_clause[5][43] 	= 1'b1;
			partial_clause[5][44] 	= 1'b1;
			partial_clause[5][45] 	= 1'b0;
			partial_clause[5][46] 	= 1'b1;
			partial_clause[5][47] 	= 1'b1;
			partial_clause[5][48] 	= 1'b1;
			partial_clause[5][49] 	= 1'b1;
			partial_clause[5][50] 	= 1'b1;
			partial_clause[5][51] 	= 1'b1;
			partial_clause[5][52] 	= 1'b0;
			partial_clause[5][53] 	= 1'b1;
			partial_clause[5][54] 	= 1'b1;
			partial_clause[5][55] 	= 1'b1;
			partial_clause[5][56] 	= 1'b1;
			partial_clause[5][57] 	= x[24];
			partial_clause[5][58] 	= 1'b1;
			partial_clause[5][59] 	= 1'b1;
			partial_clause[5][60] 	= 1'b1;
			partial_clause[5][61] 	= 1'b0;
			partial_clause[5][62] 	= 1'b1;
			partial_clause[5][63] 	= 1'b1;
			partial_clause[5][64] 	= 1'b1;
			partial_clause[5][65] 	= 1'b1;
			partial_clause[5][66] 	= 1'b1;
			partial_clause[5][67] 	= 1'b1;
			partial_clause[5][68] 	= 1'b1;
			partial_clause[5][69] 	= 1'b1;
			partial_clause[5][70] 	= 1'b0;
			partial_clause[5][71] 	= 1'b1;
			partial_clause[5][72] 	= x[10];
			partial_clause[5][73] 	= 1'b1;
			partial_clause[5][74] 	= 1'b1;
			partial_clause[5][75] 	= 1'b1;
			partial_clause[5][76] 	= 1'b1;
			partial_clause[5][77] 	= x[15];
			partial_clause[5][78] 	= 1'b1;
			partial_clause[5][79] 	= 1'b1;
			partial_clause[5][80] 	= 1'b1;
			partial_clause[5][81] 	= 1'b1;
			partial_clause[5][82] 	= 1'b1;
			partial_clause[5][83] 	= 1'b1;
			partial_clause[5][84] 	= 1'b1;
			partial_clause[5][85] 	= 1'b1;
			partial_clause[5][86] 	= x[27];
			partial_clause[5][87] 	= 1'b1;
			partial_clause[5][88] 	= 1'b1;
			partial_clause[5][89] 	= 1'b1;
			partial_clause[5][90] 	= 1'b1;
			partial_clause[5][91] 	= 1'b1;
			partial_clause[5][92] 	= 1'b1;
			partial_clause[5][93] 	= 1'b0;
			partial_clause[5][94] 	= 1'b1;
			partial_clause[5][95] 	= 1'b1;
			partial_clause[5][96] 	= 1'b1;
			partial_clause[5][97] 	= 1'b1;
			partial_clause[5][98] 	= 1'b1;
			partial_clause[5][99] 	= 1'b1;
			partial_clause[5][100] 	= 1'b1;
			partial_clause[5][101] 	= 1'b1;
			partial_clause[5][102] 	= 1'b0;
			partial_clause[5][103] 	= 1'b1;
			partial_clause[5][104] 	= 1'b1;
			partial_clause[5][105] 	= 1'b1;
			partial_clause[5][106] 	= 1'b1;
			partial_clause[5][107] 	= 1'b1;
			partial_clause[5][108] 	= 1'b1;
			partial_clause[5][109] 	= 1'b1;
			partial_clause[5][110] 	= 1'b1;
			partial_clause[5][111] 	= 1'b1;
			partial_clause[5][112] 	= 1'b1;
			partial_clause[5][113] 	= 1'b1;
			partial_clause[5][114] 	= 1'b1;
			partial_clause[5][115] 	= 1'b1;
			partial_clause[5][116] 	= 1'b1;
			partial_clause[5][117] 	= 1'b1;
			partial_clause[5][118] 	= 1'b0;
			partial_clause[5][119] 	= 1'b1;
			partial_clause[5][120] 	= 1'b1;
			partial_clause[5][121] 	= 1'b1;
			partial_clause[5][122] 	= 1'b1;
			partial_clause[5][123] 	= 1'b1;
			partial_clause[5][124] 	= 1'b1;
			partial_clause[5][125] 	= 1'b1;
			partial_clause[5][126] 	= 1'b0;
			partial_clause[5][127] 	= 1'b1;
			partial_clause[5][128] 	= 1'b1;
			partial_clause[5][129] 	= 1'b1;
			partial_clause[5][130] 	= 1'b1;
			partial_clause[5][131] 	= 1'b1;
			partial_clause[5][132] 	= 1'b1;
			partial_clause[5][133] 	= 1'b1;
			partial_clause[5][134] 	= 1'b1;
			partial_clause[5][135] 	= 1'b1;
			partial_clause[5][136] 	= 1'b1;
			partial_clause[5][137] 	= 1'b1;
			partial_clause[5][138] 	= 1'b1;
			partial_clause[5][139] 	= 1'b1;
			partial_clause[5][140] 	= 1'b1;
			partial_clause[5][141] 	= 1'b1;
			partial_clause[5][142] 	= 1'b1;
			partial_clause[5][143] 	= 1'b1;
			partial_clause[5][144] 	= 1'b1;
			partial_clause[5][145] 	= 1'b1;
			partial_clause[5][146] 	= 1'b1;
			partial_clause[5][147] 	= 1'b1;
			partial_clause[5][148] 	= 1'b1;
			partial_clause[5][149] 	= 1'b1;
			partial_clause[5][150] 	= 1'b1;
			partial_clause[5][151] 	= 1'b1;
			partial_clause[5][152] 	= 1'b1;
			partial_clause[5][153] 	= x[27];
			partial_clause[5][154] 	= 1'b1;
			partial_clause[5][155] 	= 1'b1;
			partial_clause[5][156] 	= 1'b1;
			partial_clause[5][157] 	= 1'b1;
			partial_clause[5][158] 	= 1'b1;
			partial_clause[5][159] 	= 1'b1;
			partial_clause[5][160] 	= 1'b1;
			partial_clause[5][161] 	= 1'b1;
			partial_clause[5][162] 	= 1'b1;
			partial_clause[5][163] 	= 1'b1;
			partial_clause[5][164] 	= 1'b1;
			partial_clause[5][165] 	= 1'b1;
			partial_clause[5][166] 	= 1'b1;
			partial_clause[5][167] 	= 1'b1;
			partial_clause[5][168] 	= 1'b1;
			partial_clause[5][169] 	= 1'b1;
			partial_clause[5][170] 	= 1'b1;
			partial_clause[5][171] 	= 1'b1;
			partial_clause[5][172] 	= 1'b1;
			partial_clause[5][173] 	= 1'b0;
			partial_clause[5][174] 	= 1'b1;
			partial_clause[5][175] 	= 1'b1;
			partial_clause[5][176] 	= 1'b1;
			partial_clause[5][177] 	= 1'b1;
			partial_clause[5][178] 	= 1'b1;
			partial_clause[5][179] 	= 1'b1;
			partial_clause[5][180] 	= 1'b1;
			partial_clause[5][181] 	= 1'b1;
			partial_clause[5][182] 	= 1'b1;
			partial_clause[5][183] 	= 1'b1;
			partial_clause[5][184] 	= 1'b1;
			partial_clause[5][185] 	= 1'b1;
			partial_clause[5][186] 	= 1'b1;
			partial_clause[5][187] 	= 1'b1;
			partial_clause[5][188] 	= 1'b1;
			partial_clause[5][189] 	= 1'b1;
			partial_clause[5][190] 	= 1'b1;
			partial_clause[5][191] 	= 1'b1;
			partial_clause[5][192] 	= 1'b1;
			partial_clause[5][193] 	= 1'b1;
			partial_clause[5][194] 	= 1'b1;
			partial_clause[5][195] 	= 1'b0;
			partial_clause[5][196] 	= 1'b1;
			partial_clause[5][197] 	= 1'b0;
			partial_clause[5][198] 	= 1'b1;
			partial_clause[5][199] 	= 1'b1;
			// Class 6
			partial_clause[6][0] 	= 1'b1;
			partial_clause[6][1] 	= 1'b1;
			partial_clause[6][2] 	= 1'b1;
			partial_clause[6][3] 	= 1'b1;
			partial_clause[6][4] 	= 1'b1;
			partial_clause[6][5] 	= x[60];
			partial_clause[6][6] 	= 1'b1;
			partial_clause[6][7] 	= x[33];
			partial_clause[6][8] 	= 1'b0;
			partial_clause[6][9] 	= 1'b1;
			partial_clause[6][10] 	= 1'b1;
			partial_clause[6][11] 	= 1'b1;
			partial_clause[6][12] 	= x[31];
			partial_clause[6][13] 	= x[11];
			partial_clause[6][14] 	= 1'b1;
			partial_clause[6][15] 	= 1'b1;
			partial_clause[6][16] 	= 1'b1;
			partial_clause[6][17] 	= 1'b1;
			partial_clause[6][18] 	= x[23];
			partial_clause[6][19] 	= 1'b1;
			partial_clause[6][20] 	= 1'b1;
			partial_clause[6][21] 	= 1'b1;
			partial_clause[6][22] 	= 1'b1;
			partial_clause[6][23] 	= 1'b1;
			partial_clause[6][24] 	= 1'b1;
			partial_clause[6][25] 	= 1'b1;
			partial_clause[6][26] 	= 1'b0;
			partial_clause[6][27] 	= x[34];
			partial_clause[6][28] 	= 1'b1;
			partial_clause[6][29] 	= 1'b1;
			partial_clause[6][30] 	= 1'b1;
			partial_clause[6][31] 	= 1'b1;
			partial_clause[6][32] 	= 1'b0;
			partial_clause[6][33] 	= x[54];
			partial_clause[6][34] 	= 1'b0;
			partial_clause[6][35] 	= x[63];
			partial_clause[6][36] 	= 1'b1;
			partial_clause[6][37] 	= 1'b1;
			partial_clause[6][38] 	= 1'b1;
			partial_clause[6][39] 	= x[20];
			partial_clause[6][40] 	= 1'b1;
			partial_clause[6][41] 	= 1'b1;
			partial_clause[6][42] 	= 1'b1;
			partial_clause[6][43] 	= 1'b1;
			partial_clause[6][44] 	= 1'b1;
			partial_clause[6][45] 	= 1'b1;
			partial_clause[6][46] 	= 1'b1;
			partial_clause[6][47] 	= 1'b1;
			partial_clause[6][48] 	= 1'b1;
			partial_clause[6][49] 	= 1'b1;
			partial_clause[6][50] 	= 1'b1;
			partial_clause[6][51] 	= 1'b1;
			partial_clause[6][52] 	= 1'b1;
			partial_clause[6][53] 	= 1'b1;
			partial_clause[6][54] 	= 1'b1;
			partial_clause[6][55] 	= 1'b1;
			partial_clause[6][56] 	= 1'b1;
			partial_clause[6][57] 	= x[32];
			partial_clause[6][58] 	= 1'b1;
			partial_clause[6][59] 	= 1'b0;
			partial_clause[6][60] 	= 1'b1;
			partial_clause[6][61] 	= 1'b1;
			partial_clause[6][62] 	= 1'b1;
			partial_clause[6][63] 	= 1'b1;
			partial_clause[6][64] 	= 1'b1;
			partial_clause[6][65] 	= 1'b0;
			partial_clause[6][66] 	= 1'b1;
			partial_clause[6][67] 	= 1'b1;
			partial_clause[6][68] 	= 1'b1;
			partial_clause[6][69] 	= 1'b1;
			partial_clause[6][70] 	= 1'b0;
			partial_clause[6][71] 	= 1'b1;
			partial_clause[6][72] 	= 1'b1;
			partial_clause[6][73] 	= 1'b1;
			partial_clause[6][74] 	= 1'b1;
			partial_clause[6][75] 	= 1'b1;
			partial_clause[6][76] 	= 1'b1;
			partial_clause[6][77] 	= 1'b0;
			partial_clause[6][78] 	= 1'b1;
			partial_clause[6][79] 	= 1'b1;
			partial_clause[6][80] 	= x[11];
			partial_clause[6][81] 	= 1'b0;
			partial_clause[6][82] 	= 1'b1;
			partial_clause[6][83] 	= 1'b0;
			partial_clause[6][84] 	= 1'b1;
			partial_clause[6][85] 	= 1'b1;
			partial_clause[6][86] 	= x[5];
			partial_clause[6][87] 	= x[28];
			partial_clause[6][88] 	= 1'b1;
			partial_clause[6][89] 	= 1'b1;
			partial_clause[6][90] 	= 1'b1;
			partial_clause[6][91] 	= 1'b1;
			partial_clause[6][92] 	= x[25];
			partial_clause[6][93] 	= 1'b1;
			partial_clause[6][94] 	= 1'b1;
			partial_clause[6][95] 	= 1'b1;
			partial_clause[6][96] 	= 1'b1;
			partial_clause[6][97] 	= 1'b1;
			partial_clause[6][98] 	= 1'b1;
			partial_clause[6][99] 	= 1'b1;
			partial_clause[6][100] 	= 1'b1;
			partial_clause[6][101] 	= 1'b1;
			partial_clause[6][102] 	= 1'b1;
			partial_clause[6][103] 	= 1'b0;
			partial_clause[6][104] 	= 1'b1;
			partial_clause[6][105] 	= 1'b1;
			partial_clause[6][106] 	= 1'b1;
			partial_clause[6][107] 	= 1'b1;
			partial_clause[6][108] 	= 1'b1;
			partial_clause[6][109] 	= 1'b0;
			partial_clause[6][110] 	= 1'b1;
			partial_clause[6][111] 	= 1'b1;
			partial_clause[6][112] 	= 1'b1;
			partial_clause[6][113] 	= 1'b1;
			partial_clause[6][114] 	= 1'b1;
			partial_clause[6][115] 	= 1'b1;
			partial_clause[6][116] 	= 1'b1;
			partial_clause[6][117] 	= 1'b1;
			partial_clause[6][118] 	= 1'b1;
			partial_clause[6][119] 	= 1'b1;
			partial_clause[6][120] 	= ~x[44];
			partial_clause[6][121] 	= 1'b1;
			partial_clause[6][122] 	= 1'b1;
			partial_clause[6][123] 	= 1'b1;
			partial_clause[6][124] 	= 1'b1;
			partial_clause[6][125] 	= ~x[61];
			partial_clause[6][126] 	= 1'b1;
			partial_clause[6][127] 	= 1'b1;
			partial_clause[6][128] 	= 1'b1;
			partial_clause[6][129] 	= 1'b1;
			partial_clause[6][130] 	= 1'b1;
			partial_clause[6][131] 	= 1'b1;
			partial_clause[6][132] 	= 1'b1;
			partial_clause[6][133] 	= 1'b1;
			partial_clause[6][134] 	= 1'b1;
			partial_clause[6][135] 	= 1'b1;
			partial_clause[6][136] 	= 1'b1;
			partial_clause[6][137] 	= 1'b1;
			partial_clause[6][138] 	= 1'b1;
			partial_clause[6][139] 	= 1'b1;
			partial_clause[6][140] 	= 1'b1;
			partial_clause[6][141] 	= 1'b1;
			partial_clause[6][142] 	= 1'b1;
			partial_clause[6][143] 	= 1'b1;
			partial_clause[6][144] 	= 1'b1;
			partial_clause[6][145] 	= 1'b0;
			partial_clause[6][146] 	= 1'b1;
			partial_clause[6][147] 	= 1'b1;
			partial_clause[6][148] 	= 1'b1;
			partial_clause[6][149] 	= 1'b1;
			partial_clause[6][150] 	= 1'b1;
			partial_clause[6][151] 	= 1'b1;
			partial_clause[6][152] 	= 1'b1;
			partial_clause[6][153] 	= 1'b1;
			partial_clause[6][154] 	= 1'b1;
			partial_clause[6][155] 	= 1'b1;
			partial_clause[6][156] 	= 1'b1;
			partial_clause[6][157] 	= 1'b1;
			partial_clause[6][158] 	= 1'b1;
			partial_clause[6][159] 	= 1'b1;
			partial_clause[6][160] 	= 1'b1;
			partial_clause[6][161] 	= 1'b1;
			partial_clause[6][162] 	= 1'b1;
			partial_clause[6][163] 	= 1'b1;
			partial_clause[6][164] 	= 1'b1;
			partial_clause[6][165] 	= 1'b1;
			partial_clause[6][166] 	= 1'b1;
			partial_clause[6][167] 	= 1'b1;
			partial_clause[6][168] 	= 1'b1;
			partial_clause[6][169] 	= 1'b1;
			partial_clause[6][170] 	= 1'b1;
			partial_clause[6][171] 	= 1'b1;
			partial_clause[6][172] 	= 1'b1;
			partial_clause[6][173] 	= 1'b1;
			partial_clause[6][174] 	= 1'b1;
			partial_clause[6][175] 	= 1'b1;
			partial_clause[6][176] 	= 1'b1;
			partial_clause[6][177] 	= 1'b1;
			partial_clause[6][178] 	= 1'b1;
			partial_clause[6][179] 	= 1'b1;
			partial_clause[6][180] 	= 1'b1;
			partial_clause[6][181] 	= 1'b1;
			partial_clause[6][182] 	= 1'b1;
			partial_clause[6][183] 	= 1'b1;
			partial_clause[6][184] 	= 1'b1;
			partial_clause[6][185] 	= 1'b1;
			partial_clause[6][186] 	= 1'b1;
			partial_clause[6][187] 	= 1'b1;
			partial_clause[6][188] 	= 1'b1;
			partial_clause[6][189] 	= 1'b1;
			partial_clause[6][190] 	= 1'b1;
			partial_clause[6][191] 	= 1'b1;
			partial_clause[6][192] 	= 1'b1;
			partial_clause[6][193] 	= 1'b1;
			partial_clause[6][194] 	= 1'b1;
			partial_clause[6][195] 	= 1'b1;
			partial_clause[6][196] 	= 1'b1;
			partial_clause[6][197] 	= 1'b1;
			partial_clause[6][198] 	= 1'b1;
			partial_clause[6][199] 	= 1'b1;
			// Class 7
			partial_clause[7][0] 	= 1'b1;
			partial_clause[7][1] 	= 1'b1;
			partial_clause[7][2] 	= 1'b1;
			partial_clause[7][3] 	= x[17];
			partial_clause[7][4] 	= 1'b1;
			partial_clause[7][5] 	= 1'b1;
			partial_clause[7][6] 	= 1'b1;
			partial_clause[7][7] 	= 1'b0;
			partial_clause[7][8] 	= 1'b1;
			partial_clause[7][9] 	= 1'b1;
			partial_clause[7][10] 	= 1'b1;
			partial_clause[7][11] 	= 1'b1;
			partial_clause[7][12] 	= 1'b0;
			partial_clause[7][13] 	= x[56];
			partial_clause[7][14] 	= 1'b1;
			partial_clause[7][15] 	= 1'b1;
			partial_clause[7][16] 	= 1'b1;
			partial_clause[7][17] 	= 1'b1;
			partial_clause[7][18] 	= 1'b1;
			partial_clause[7][19] 	= 1'b1;
			partial_clause[7][20] 	= 1'b1;
			partial_clause[7][21] 	= 1'b1;
			partial_clause[7][22] 	= 1'b1;
			partial_clause[7][23] 	= 1'b1;
			partial_clause[7][24] 	= 1'b1;
			partial_clause[7][25] 	= 1'b1;
			partial_clause[7][26] 	= 1'b1;
			partial_clause[7][27] 	= x[8];
			partial_clause[7][28] 	= 1'b1;
			partial_clause[7][29] 	= x[51];
			partial_clause[7][30] 	= 1'b1;
			partial_clause[7][31] 	= 1'b1;
			partial_clause[7][32] 	= 1'b0;
			partial_clause[7][33] 	= 1'b1;
			partial_clause[7][34] 	= 1'b1;
			partial_clause[7][35] 	= x[48];
			partial_clause[7][36] 	= 1'b1;
			partial_clause[7][37] 	= 1'b1;
			partial_clause[7][38] 	= 1'b1;
			partial_clause[7][39] 	= 1'b1;
			partial_clause[7][40] 	= 1'b1;
			partial_clause[7][41] 	= 1'b1;
			partial_clause[7][42] 	= 1'b1;
			partial_clause[7][43] 	= 1'b1;
			partial_clause[7][44] 	= 1'b1;
			partial_clause[7][45] 	= 1'b1;
			partial_clause[7][46] 	= 1'b0;
			partial_clause[7][47] 	= 1'b1;
			partial_clause[7][48] 	= 1'b1;
			partial_clause[7][49] 	= 1'b0;
			partial_clause[7][50] 	= 1'b1;
			partial_clause[7][51] 	= 1'b1;
			partial_clause[7][52] 	= 1'b0;
			partial_clause[7][53] 	= 1'b1;
			partial_clause[7][54] 	= 1'b0;
			partial_clause[7][55] 	= x[48];
			partial_clause[7][56] 	= 1'b0;
			partial_clause[7][57] 	= 1'b1;
			partial_clause[7][58] 	= 1'b1;
			partial_clause[7][59] 	= x[6];
			partial_clause[7][60] 	= 1'b1;
			partial_clause[7][61] 	= 1'b1;
			partial_clause[7][62] 	= 1'b1;
			partial_clause[7][63] 	= 1'b1;
			partial_clause[7][64] 	= 1'b1;
			partial_clause[7][65] 	= 1'b1;
			partial_clause[7][66] 	= 1'b1;
			partial_clause[7][67] 	= 1'b1;
			partial_clause[7][68] 	= 1'b1;
			partial_clause[7][69] 	= 1'b1;
			partial_clause[7][70] 	= 1'b1;
			partial_clause[7][71] 	= 1'b1;
			partial_clause[7][72] 	= 1'b1;
			partial_clause[7][73] 	= 1'b1;
			partial_clause[7][74] 	= 1'b1;
			partial_clause[7][75] 	= 1'b1;
			partial_clause[7][76] 	= 1'b1;
			partial_clause[7][77] 	= 1'b1;
			partial_clause[7][78] 	= 1'b1;
			partial_clause[7][79] 	= 1'b0;
			partial_clause[7][80] 	= 1'b0;
			partial_clause[7][81] 	= 1'b1;
			partial_clause[7][82] 	= 1'b1;
			partial_clause[7][83] 	= 1'b1;
			partial_clause[7][84] 	= 1'b1;
			partial_clause[7][85] 	= x[53];
			partial_clause[7][86] 	= 1'b1;
			partial_clause[7][87] 	= 1'b1;
			partial_clause[7][88] 	= x[24];
			partial_clause[7][89] 	= 1'b1;
			partial_clause[7][90] 	= 1'b1;
			partial_clause[7][91] 	= 1'b1;
			partial_clause[7][92] 	= 1'b1;
			partial_clause[7][93] 	= 1'b1;
			partial_clause[7][94] 	= x[10];
			partial_clause[7][95] 	= 1'b1;
			partial_clause[7][96] 	= 1'b1;
			partial_clause[7][97] 	= 1'b1;
			partial_clause[7][98] 	= 1'b1;
			partial_clause[7][99] 	= 1'b1;
			partial_clause[7][100] 	= 1'b1;
			partial_clause[7][101] 	= 1'b1;
			partial_clause[7][102] 	= 1'b1;
			partial_clause[7][103] 	= 1'b1;
			partial_clause[7][104] 	= 1'b1;
			partial_clause[7][105] 	= 1'b1;
			partial_clause[7][106] 	= 1'b1;
			partial_clause[7][107] 	= 1'b1;
			partial_clause[7][108] 	= 1'b1;
			partial_clause[7][109] 	= 1'b1;
			partial_clause[7][110] 	= 1'b1;
			partial_clause[7][111] 	= 1'b1;
			partial_clause[7][112] 	= 1'b1;
			partial_clause[7][113] 	= 1'b1;
			partial_clause[7][114] 	= 1'b1;
			partial_clause[7][115] 	= 1'b1;
			partial_clause[7][116] 	= 1'b1;
			partial_clause[7][117] 	= 1'b1;
			partial_clause[7][118] 	= 1'b1;
			partial_clause[7][119] 	= 1'b1;
			partial_clause[7][120] 	= 1'b0;
			partial_clause[7][121] 	= 1'b0;
			partial_clause[7][122] 	= 1'b1;
			partial_clause[7][123] 	= 1'b1;
			partial_clause[7][124] 	= 1'b1;
			partial_clause[7][125] 	= 1'b1;
			partial_clause[7][126] 	= 1'b1;
			partial_clause[7][127] 	= 1'b0;
			partial_clause[7][128] 	= 1'b1;
			partial_clause[7][129] 	= 1'b1;
			partial_clause[7][130] 	= 1'b1;
			partial_clause[7][131] 	= 1'b1;
			partial_clause[7][132] 	= 1'b1;
			partial_clause[7][133] 	= 1'b1;
			partial_clause[7][134] 	= 1'b1;
			partial_clause[7][135] 	= 1'b1;
			partial_clause[7][136] 	= 1'b1;
			partial_clause[7][137] 	= 1'b1;
			partial_clause[7][138] 	= 1'b1;
			partial_clause[7][139] 	= 1'b1;
			partial_clause[7][140] 	= 1'b1;
			partial_clause[7][141] 	= 1'b1;
			partial_clause[7][142] 	= 1'b1;
			partial_clause[7][143] 	= 1'b1;
			partial_clause[7][144] 	= 1'b1;
			partial_clause[7][145] 	= 1'b1;
			partial_clause[7][146] 	= 1'b1;
			partial_clause[7][147] 	= 1'b1;
			partial_clause[7][148] 	= 1'b1;
			partial_clause[7][149] 	= 1'b1;
			partial_clause[7][150] 	= 1'b1;
			partial_clause[7][151] 	= 1'b1;
			partial_clause[7][152] 	= 1'b1;
			partial_clause[7][153] 	= 1'b1;
			partial_clause[7][154] 	= 1'b1;
			partial_clause[7][155] 	= 1'b1;
			partial_clause[7][156] 	= 1'b1;
			partial_clause[7][157] 	= 1'b1;
			partial_clause[7][158] 	= 1'b1;
			partial_clause[7][159] 	= 1'b1;
			partial_clause[7][160] 	= 1'b1;
			partial_clause[7][161] 	= 1'b1;
			partial_clause[7][162] 	= 1'b1;
			partial_clause[7][163] 	= 1'b1;
			partial_clause[7][164] 	= 1'b1;
			partial_clause[7][165] 	= 1'b1;
			partial_clause[7][166] 	= 1'b1;
			partial_clause[7][167] 	= 1'b1;
			partial_clause[7][168] 	= 1'b1;
			partial_clause[7][169] 	= 1'b0;
			partial_clause[7][170] 	= 1'b1;
			partial_clause[7][171] 	= 1'b1;
			partial_clause[7][172] 	= 1'b1;
			partial_clause[7][173] 	= 1'b1;
			partial_clause[7][174] 	= 1'b1;
			partial_clause[7][175] 	= 1'b1;
			partial_clause[7][176] 	= 1'b1;
			partial_clause[7][177] 	= 1'b1;
			partial_clause[7][178] 	= 1'b1;
			partial_clause[7][179] 	= 1'b1;
			partial_clause[7][180] 	= 1'b1;
			partial_clause[7][181] 	= 1'b1;
			partial_clause[7][182] 	= 1'b1;
			partial_clause[7][183] 	= 1'b0;
			partial_clause[7][184] 	= 1'b1;
			partial_clause[7][185] 	= 1'b1;
			partial_clause[7][186] 	= 1'b1;
			partial_clause[7][187] 	= 1'b1;
			partial_clause[7][188] 	= 1'b1;
			partial_clause[7][189] 	= 1'b1;
			partial_clause[7][190] 	= 1'b1;
			partial_clause[7][191] 	= 1'b1;
			partial_clause[7][192] 	= 1'b1;
			partial_clause[7][193] 	= 1'b1;
			partial_clause[7][194] 	= 1'b1;
			partial_clause[7][195] 	= 1'b0;
			partial_clause[7][196] 	= 1'b1;
			partial_clause[7][197] 	= 1'b1;
			partial_clause[7][198] 	= 1'b1;
			partial_clause[7][199] 	= 1'b1;
			// Class 8
			partial_clause[8][0] 	= 1'b1;
			partial_clause[8][1] 	= 1'b1;
			partial_clause[8][2] 	= 1'b1;
			partial_clause[8][3] 	= 1'b0;
			partial_clause[8][4] 	= 1'b1;
			partial_clause[8][5] 	= 1'b1;
			partial_clause[8][6] 	= 1'b1;
			partial_clause[8][7] 	= x[52];
			partial_clause[8][8] 	= 1'b1;
			partial_clause[8][9] 	= 1'b1;
			partial_clause[8][10] 	= 1'b1;
			partial_clause[8][11] 	= 1'b1;
			partial_clause[8][12] 	= 1'b1;
			partial_clause[8][13] 	= 1'b1;
			partial_clause[8][14] 	= 1'b1;
			partial_clause[8][15] 	= 1'b1;
			partial_clause[8][16] 	= ~x[23];
			partial_clause[8][17] 	= 1'b1;
			partial_clause[8][18] 	= 1'b1;
			partial_clause[8][19] 	= 1'b1;
			partial_clause[8][20] 	= x[25];
			partial_clause[8][21] 	= 1'b1;
			partial_clause[8][22] 	= 1'b1;
			partial_clause[8][23] 	= 1'b1;
			partial_clause[8][24] 	= 1'b1;
			partial_clause[8][25] 	= 1'b1;
			partial_clause[8][26] 	= 1'b1;
			partial_clause[8][27] 	= 1'b1;
			partial_clause[8][28] 	= 1'b1;
			partial_clause[8][29] 	= 1'b1;
			partial_clause[8][30] 	= 1'b1;
			partial_clause[8][31] 	= 1'b1;
			partial_clause[8][32] 	= 1'b1;
			partial_clause[8][33] 	= 1'b1;
			partial_clause[8][34] 	= 1'b1;
			partial_clause[8][35] 	= 1'b1;
			partial_clause[8][36] 	= 1'b1;
			partial_clause[8][37] 	= 1'b1;
			partial_clause[8][38] 	= 1'b1;
			partial_clause[8][39] 	= 1'b1;
			partial_clause[8][40] 	= x[36];
			partial_clause[8][41] 	= 1'b1;
			partial_clause[8][42] 	= 1'b1;
			partial_clause[8][43] 	= 1'b1;
			partial_clause[8][44] 	= 1'b1;
			partial_clause[8][45] 	= 1'b1;
			partial_clause[8][46] 	= 1'b1;
			partial_clause[8][47] 	= 1'b1;
			partial_clause[8][48] 	= 1'b1;
			partial_clause[8][49] 	= 1'b0;
			partial_clause[8][50] 	= 1'b1;
			partial_clause[8][51] 	= 1'b1;
			partial_clause[8][52] 	= 1'b1;
			partial_clause[8][53] 	= 1'b1;
			partial_clause[8][54] 	= 1'b1;
			partial_clause[8][55] 	= 1'b1;
			partial_clause[8][56] 	= 1'b1;
			partial_clause[8][57] 	= 1'b1;
			partial_clause[8][58] 	= 1'b1;
			partial_clause[8][59] 	= 1'b1;
			partial_clause[8][60] 	= 1'b1;
			partial_clause[8][61] 	= 1'b1;
			partial_clause[8][62] 	= 1'b1;
			partial_clause[8][63] 	= 1'b1;
			partial_clause[8][64] 	= 1'b1;
			partial_clause[8][65] 	= 1'b1;
			partial_clause[8][66] 	= 1'b1;
			partial_clause[8][67] 	= 1'b1;
			partial_clause[8][68] 	= 1'b1;
			partial_clause[8][69] 	= 1'b1;
			partial_clause[8][70] 	= 1'b1;
			partial_clause[8][71] 	= 1'b1;
			partial_clause[8][72] 	= 1'b1;
			partial_clause[8][73] 	= 1'b1;
			partial_clause[8][74] 	= 1'b1;
			partial_clause[8][75] 	= 1'b1;
			partial_clause[8][76] 	= 1'b1;
			partial_clause[8][77] 	= 1'b1;
			partial_clause[8][78] 	= 1'b1;
			partial_clause[8][79] 	= 1'b1;
			partial_clause[8][80] 	= 1'b1;
			partial_clause[8][81] 	= 1'b1;
			partial_clause[8][82] 	= 1'b1;
			partial_clause[8][83] 	= 1'b1;
			partial_clause[8][84] 	= 1'b1;
			partial_clause[8][85] 	= 1'b1;
			partial_clause[8][86] 	= 1'b1;
			partial_clause[8][87] 	= 1'b1;
			partial_clause[8][88] 	= 1'b0;
			partial_clause[8][89] 	= 1'b1;
			partial_clause[8][90] 	= 1'b1;
			partial_clause[8][91] 	= 1'b1;
			partial_clause[8][92] 	= 1'b1;
			partial_clause[8][93] 	= 1'b1;
			partial_clause[8][94] 	= 1'b1;
			partial_clause[8][95] 	= 1'b1;
			partial_clause[8][96] 	= 1'b0;
			partial_clause[8][97] 	= 1'b1;
			partial_clause[8][98] 	= 1'b1;
			partial_clause[8][99] 	= 1'b1;
			partial_clause[8][100] 	= 1'b1;
			partial_clause[8][101] 	= 1'b0;
			partial_clause[8][102] 	= 1'b1;
			partial_clause[8][103] 	= 1'b1;
			partial_clause[8][104] 	= 1'b1;
			partial_clause[8][105] 	= 1'b1;
			partial_clause[8][106] 	= 1'b1;
			partial_clause[8][107] 	= 1'b1;
			partial_clause[8][108] 	= 1'b1;
			partial_clause[8][109] 	= 1'b1;
			partial_clause[8][110] 	= 1'b1;
			partial_clause[8][111] 	= 1'b1;
			partial_clause[8][112] 	= 1'b1;
			partial_clause[8][113] 	= 1'b1;
			partial_clause[8][114] 	= ~x[44];
			partial_clause[8][115] 	= 1'b1;
			partial_clause[8][116] 	= 1'b1;
			partial_clause[8][117] 	= 1'b1;
			partial_clause[8][118] 	= 1'b1;
			partial_clause[8][119] 	= 1'b1;
			partial_clause[8][120] 	= 1'b1;
			partial_clause[8][121] 	= 1'b1;
			partial_clause[8][122] 	= 1'b1;
			partial_clause[8][123] 	= 1'b1;
			partial_clause[8][124] 	= 1'b0;
			partial_clause[8][125] 	= 1'b1;
			partial_clause[8][126] 	= 1'b1;
			partial_clause[8][127] 	= ~x[1];
			partial_clause[8][128] 	= 1'b1;
			partial_clause[8][129] 	= 1'b1;
			partial_clause[8][130] 	= 1'b1;
			partial_clause[8][131] 	= 1'b1;
			partial_clause[8][132] 	= 1'b1;
			partial_clause[8][133] 	= 1'b1;
			partial_clause[8][134] 	= 1'b1;
			partial_clause[8][135] 	= 1'b1;
			partial_clause[8][136] 	= x[37];
			partial_clause[8][137] 	= 1'b1;
			partial_clause[8][138] 	= 1'b1;
			partial_clause[8][139] 	= 1'b1;
			partial_clause[8][140] 	= 1'b1;
			partial_clause[8][141] 	= ~x[38];
			partial_clause[8][142] 	= x[19];
			partial_clause[8][143] 	= 1'b1;
			partial_clause[8][144] 	= 1'b1;
			partial_clause[8][145] 	= 1'b1;
			partial_clause[8][146] 	= x[56];
			partial_clause[8][147] 	= 1'b1;
			partial_clause[8][148] 	= 1'b1;
			partial_clause[8][149] 	= x[27];
			partial_clause[8][150] 	= 1'b1;
			partial_clause[8][151] 	= 1'b1;
			partial_clause[8][152] 	= 1'b1;
			partial_clause[8][153] 	= ~x[42];
			partial_clause[8][154] 	= 1'b1;
			partial_clause[8][155] 	= 1'b1;
			partial_clause[8][156] 	= 1'b1;
			partial_clause[8][157] 	= 1'b1;
			partial_clause[8][158] 	= 1'b1;
			partial_clause[8][159] 	= 1'b0;
			partial_clause[8][160] 	= 1'b1;
			partial_clause[8][161] 	= 1'b1;
			partial_clause[8][162] 	= 1'b1;
			partial_clause[8][163] 	= ~x[27];
			partial_clause[8][164] 	= 1'b1;
			partial_clause[8][165] 	= 1'b1;
			partial_clause[8][166] 	= 1'b1;
			partial_clause[8][167] 	= 1'b1;
			partial_clause[8][168] 	= 1'b1;
			partial_clause[8][169] 	= 1'b1;
			partial_clause[8][170] 	= 1'b1;
			partial_clause[8][171] 	= 1'b1;
			partial_clause[8][172] 	= 1'b1;
			partial_clause[8][173] 	= 1'b1;
			partial_clause[8][174] 	= 1'b1;
			partial_clause[8][175] 	= 1'b1;
			partial_clause[8][176] 	= 1'b1;
			partial_clause[8][177] 	= 1'b1;
			partial_clause[8][178] 	= 1'b1;
			partial_clause[8][179] 	= 1'b1;
			partial_clause[8][180] 	= 1'b1;
			partial_clause[8][181] 	= 1'b0;
			partial_clause[8][182] 	= 1'b1;
			partial_clause[8][183] 	= ~x[40];
			partial_clause[8][184] 	= 1'b1;
			partial_clause[8][185] 	= 1'b1;
			partial_clause[8][186] 	= 1'b1;
			partial_clause[8][187] 	= 1'b1;
			partial_clause[8][188] 	= 1'b1;
			partial_clause[8][189] 	= 1'b0;
			partial_clause[8][190] 	= 1'b1;
			partial_clause[8][191] 	= 1'b1;
			partial_clause[8][192] 	= 1'b1;
			partial_clause[8][193] 	= 1'b1;
			partial_clause[8][194] 	= 1'b1;
			partial_clause[8][195] 	= 1'b1;
			partial_clause[8][196] 	= 1'b1;
			partial_clause[8][197] 	= 1'b1;
			partial_clause[8][198] 	= 1'b1;
			partial_clause[8][199] 	= 1'b1;
			// Class 9
			partial_clause[9][0] 	= 1'b1;
			partial_clause[9][1] 	= 1'b0;
			partial_clause[9][2] 	= 1'b1;
			partial_clause[9][3] 	= 1'b1;
			partial_clause[9][4] 	= 1'b1;
			partial_clause[9][5] 	= 1'b0;
			partial_clause[9][6] 	= 1'b1;
			partial_clause[9][7] 	= 1'b0;
			partial_clause[9][8] 	= 1'b1;
			partial_clause[9][9] 	= x[62];
			partial_clause[9][10] 	= 1'b1;
			partial_clause[9][11] 	= 1'b1;
			partial_clause[9][12] 	= 1'b0;
			partial_clause[9][13] 	= 1'b1;
			partial_clause[9][14] 	= 1'b1;
			partial_clause[9][15] 	= 1'b1;
			partial_clause[9][16] 	= 1'b1;
			partial_clause[9][17] 	= 1'b1;
			partial_clause[9][18] 	= 1'b1;
			partial_clause[9][19] 	= 1'b1;
			partial_clause[9][20] 	= 1'b1;
			partial_clause[9][21] 	= x[55];
			partial_clause[9][22] 	= 1'b1;
			partial_clause[9][23] 	= 1'b1;
			partial_clause[9][24] 	= 1'b0;
			partial_clause[9][25] 	= 1'b1;
			partial_clause[9][26] 	= x[55];
			partial_clause[9][27] 	= 1'b1;
			partial_clause[9][28] 	= 1'b1;
			partial_clause[9][29] 	= 1'b1;
			partial_clause[9][30] 	= 1'b1;
			partial_clause[9][31] 	= 1'b1;
			partial_clause[9][32] 	= 1'b0;
			partial_clause[9][33] 	= 1'b0;
			partial_clause[9][34] 	= 1'b1;
			partial_clause[9][35] 	= 1'b1;
			partial_clause[9][36] 	= 1'b1;
			partial_clause[9][37] 	= 1'b1;
			partial_clause[9][38] 	= 1'b1;
			partial_clause[9][39] 	= 1'b1;
			partial_clause[9][40] 	= 1'b1;
			partial_clause[9][41] 	= 1'b1;
			partial_clause[9][42] 	= 1'b1;
			partial_clause[9][43] 	= 1'b1;
			partial_clause[9][44] 	= 1'b1;
			partial_clause[9][45] 	= 1'b0;
			partial_clause[9][46] 	= 1'b0;
			partial_clause[9][47] 	= x[57];
			partial_clause[9][48] 	= 1'b1;
			partial_clause[9][49] 	= 1'b1;
			partial_clause[9][50] 	= 1'b1;
			partial_clause[9][51] 	= 1'b1;
			partial_clause[9][52] 	= 1'b1;
			partial_clause[9][53] 	= 1'b0;
			partial_clause[9][54] 	= 1'b1;
			partial_clause[9][55] 	= 1'b1;
			partial_clause[9][56] 	= 1'b1;
			partial_clause[9][57] 	= 1'b0;
			partial_clause[9][58] 	= 1'b1;
			partial_clause[9][59] 	= 1'b1;
			partial_clause[9][60] 	= 1'b1;
			partial_clause[9][61] 	= 1'b1;
			partial_clause[9][62] 	= 1'b1;
			partial_clause[9][63] 	= 1'b0;
			partial_clause[9][64] 	= 1'b1;
			partial_clause[9][65] 	= 1'b1;
			partial_clause[9][66] 	= 1'b1;
			partial_clause[9][67] 	= x[40];
			partial_clause[9][68] 	= 1'b1;
			partial_clause[9][69] 	= 1'b1;
			partial_clause[9][70] 	= 1'b1;
			partial_clause[9][71] 	= 1'b1;
			partial_clause[9][72] 	= 1'b1;
			partial_clause[9][73] 	= 1'b1;
			partial_clause[9][74] 	= 1'b1;
			partial_clause[9][75] 	= 1'b1;
			partial_clause[9][76] 	= 1'b1;
			partial_clause[9][77] 	= 1'b1;
			partial_clause[9][78] 	= x[58];
			partial_clause[9][79] 	= 1'b1;
			partial_clause[9][80] 	= x[38];
			partial_clause[9][81] 	= 1'b1;
			partial_clause[9][82] 	= 1'b1;
			partial_clause[9][83] 	= x[54];
			partial_clause[9][84] 	= 1'b1;
			partial_clause[9][85] 	= 1'b1;
			partial_clause[9][86] 	= 1'b1;
			partial_clause[9][87] 	= 1'b1;
			partial_clause[9][88] 	= 1'b1;
			partial_clause[9][89] 	= 1'b1;
			partial_clause[9][90] 	= x[2];
			partial_clause[9][91] 	= 1'b1;
			partial_clause[9][92] 	= 1'b0;
			partial_clause[9][93] 	= 1'b1;
			partial_clause[9][94] 	= 1'b1;
			partial_clause[9][95] 	= 1'b1;
			partial_clause[9][96] 	= 1'b1;
			partial_clause[9][97] 	= 1'b1;
			partial_clause[9][98] 	= 1'b1;
			partial_clause[9][99] 	= 1'b1;
			partial_clause[9][100] 	= 1'b1;
			partial_clause[9][101] 	= 1'b1;
			partial_clause[9][102] 	= 1'b1;
			partial_clause[9][103] 	= 1'b1;
			partial_clause[9][104] 	= 1'b1;
			partial_clause[9][105] 	= 1'b1;
			partial_clause[9][106] 	= 1'b1;
			partial_clause[9][107] 	= 1'b1;
			partial_clause[9][108] 	= 1'b1;
			partial_clause[9][109] 	= 1'b1;
			partial_clause[9][110] 	= 1'b1;
			partial_clause[9][111] 	= 1'b1;
			partial_clause[9][112] 	= 1'b1;
			partial_clause[9][113] 	= 1'b1;
			partial_clause[9][114] 	= 1'b1;
			partial_clause[9][115] 	= 1'b1;
			partial_clause[9][116] 	= 1'b1;
			partial_clause[9][117] 	= 1'b0;
			partial_clause[9][118] 	= 1'b1;
			partial_clause[9][119] 	= 1'b1;
			partial_clause[9][120] 	= 1'b1;
			partial_clause[9][121] 	= 1'b1;
			partial_clause[9][122] 	= 1'b1;
			partial_clause[9][123] 	= 1'b1;
			partial_clause[9][124] 	= 1'b1;
			partial_clause[9][125] 	= 1'b1;
			partial_clause[9][126] 	= 1'b1;
			partial_clause[9][127] 	= 1'b1;
			partial_clause[9][128] 	= 1'b1;
			partial_clause[9][129] 	= 1'b1;
			partial_clause[9][130] 	= 1'b1;
			partial_clause[9][131] 	= 1'b1;
			partial_clause[9][132] 	= 1'b1;
			partial_clause[9][133] 	= 1'b1;
			partial_clause[9][134] 	= 1'b0;
			partial_clause[9][135] 	= 1'b0;
			partial_clause[9][136] 	= 1'b0;
			partial_clause[9][137] 	= 1'b1;
			partial_clause[9][138] 	= 1'b1;
			partial_clause[9][139] 	= 1'b1;
			partial_clause[9][140] 	= 1'b1;
			partial_clause[9][141] 	= 1'b1;
			partial_clause[9][142] 	= 1'b1;
			partial_clause[9][143] 	= 1'b1;
			partial_clause[9][144] 	= 1'b1;
			partial_clause[9][145] 	= 1'b1;
			partial_clause[9][146] 	= 1'b1;
			partial_clause[9][147] 	= 1'b1;
			partial_clause[9][148] 	= 1'b1;
			partial_clause[9][149] 	= 1'b1;
			partial_clause[9][150] 	= 1'b1;
			partial_clause[9][151] 	= 1'b1;
			partial_clause[9][152] 	= 1'b1;
			partial_clause[9][153] 	= 1'b1;
			partial_clause[9][154] 	= 1'b1;
			partial_clause[9][155] 	= 1'b1;
			partial_clause[9][156] 	= 1'b1;
			partial_clause[9][157] 	= 1'b1;
			partial_clause[9][158] 	= 1'b1;
			partial_clause[9][159] 	= 1'b1;
			partial_clause[9][160] 	= 1'b1;
			partial_clause[9][161] 	= 1'b1;
			partial_clause[9][162] 	= 1'b1;
			partial_clause[9][163] 	= 1'b1;
			partial_clause[9][164] 	= ~x[36];
			partial_clause[9][165] 	= 1'b1;
			partial_clause[9][166] 	= 1'b1;
			partial_clause[9][167] 	= 1'b1;
			partial_clause[9][168] 	= 1'b1;
			partial_clause[9][169] 	= 1'b1;
			partial_clause[9][170] 	= 1'b1;
			partial_clause[9][171] 	= 1'b1;
			partial_clause[9][172] 	= 1'b1;
			partial_clause[9][173] 	= ~x[0];
			partial_clause[9][174] 	= 1'b1;
			partial_clause[9][175] 	= 1'b1;
			partial_clause[9][176] 	= 1'b0;
			partial_clause[9][177] 	= 1'b1;
			partial_clause[9][178] 	= 1'b1;
			partial_clause[9][179] 	= 1'b1;
			partial_clause[9][180] 	= 1'b1;
			partial_clause[9][181] 	= 1'b1;
			partial_clause[9][182] 	= 1'b1;
			partial_clause[9][183] 	= 1'b1;
			partial_clause[9][184] 	= 1'b1;
			partial_clause[9][185] 	= 1'b1;
			partial_clause[9][186] 	= 1'b1;
			partial_clause[9][187] 	= 1'b1;
			partial_clause[9][188] 	= 1'b1;
			partial_clause[9][189] 	= 1'b1;
			partial_clause[9][190] 	= 1'b1;
			partial_clause[9][191] 	= 1'b1;
			partial_clause[9][192] 	= 1'b1;
			partial_clause[9][193] 	= 1'b1;
			partial_clause[9][194] 	= 1'b1;
			partial_clause[9][195] 	= 1'b1;
			partial_clause[9][196] 	= 1'b1;
			partial_clause[9][197] 	= 1'b1;
			partial_clause[9][198] 	= 1'b1;
			partial_clause[9][199] 	= 1'b1;
		end
	end
endmodule


module HCB_1 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & ~x[38];
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & ~x[3];
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & x[20];
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & x[51];
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & x[24];
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & ~x[17];
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & ~x[39];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & ~x[59];
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & ~x[39];
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			partial_clause[0][100] 	= partial_clause_prev[0][100] & 1'b1;
			partial_clause[0][101] 	= partial_clause_prev[0][101] & 1'b1;
			partial_clause[0][102] 	= partial_clause_prev[0][102] & 1'b1;
			partial_clause[0][103] 	= partial_clause_prev[0][103] & 1'b1;
			partial_clause[0][104] 	= partial_clause_prev[0][104] & 1'b1;
			partial_clause[0][105] 	= partial_clause_prev[0][105] & 1'b1;
			partial_clause[0][106] 	= partial_clause_prev[0][106] & 1'b1;
			partial_clause[0][107] 	= partial_clause_prev[0][107] & 1'b1;
			partial_clause[0][108] 	= partial_clause_prev[0][108] & 1'b1;
			partial_clause[0][109] 	= partial_clause_prev[0][109] & 1'b1;
			partial_clause[0][110] 	= partial_clause_prev[0][110] & 1'b1;
			partial_clause[0][111] 	= partial_clause_prev[0][111] & 1'b1;
			partial_clause[0][112] 	= partial_clause_prev[0][112] & 1'b1;
			partial_clause[0][113] 	= partial_clause_prev[0][113] & x[29];
			partial_clause[0][114] 	= partial_clause_prev[0][114] & 1'b1;
			partial_clause[0][115] 	= partial_clause_prev[0][115] & 1'b1;
			partial_clause[0][116] 	= partial_clause_prev[0][116] & 1'b1;
			partial_clause[0][117] 	= partial_clause_prev[0][117] & 1'b1;
			partial_clause[0][118] 	= partial_clause_prev[0][118] & 1'b1;
			partial_clause[0][119] 	= partial_clause_prev[0][119] & 1'b1;
			partial_clause[0][120] 	= partial_clause_prev[0][120] & 1'b1;
			partial_clause[0][121] 	= partial_clause_prev[0][121] & x[40];
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & 1'b1;
			partial_clause[0][124] 	= partial_clause_prev[0][124] & 1'b1;
			partial_clause[0][125] 	= partial_clause_prev[0][125] & 1'b1;
			partial_clause[0][126] 	= partial_clause_prev[0][126] & 1'b1;
			partial_clause[0][127] 	= partial_clause_prev[0][127] & 1'b1;
			partial_clause[0][128] 	= partial_clause_prev[0][128] & 1'b1;
			partial_clause[0][129] 	= partial_clause_prev[0][129] & 1'b1;
			partial_clause[0][130] 	= partial_clause_prev[0][130] & 1'b1;
			partial_clause[0][131] 	= partial_clause_prev[0][131] & 1'b1;
			partial_clause[0][132] 	= partial_clause_prev[0][132] & 1'b1;
			partial_clause[0][133] 	= partial_clause_prev[0][133] & 1'b1;
			partial_clause[0][134] 	= partial_clause_prev[0][134] & x[35];
			partial_clause[0][135] 	= partial_clause_prev[0][135] & 1'b1;
			partial_clause[0][136] 	= partial_clause_prev[0][136] & 1'b1;
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & ~x[60];
			partial_clause[0][139] 	= partial_clause_prev[0][139] & 1'b1;
			partial_clause[0][140] 	= partial_clause_prev[0][140] & 1'b1;
			partial_clause[0][141] 	= partial_clause_prev[0][141] & 1'b1;
			partial_clause[0][142] 	= partial_clause_prev[0][142] & 1'b1;
			partial_clause[0][143] 	= partial_clause_prev[0][143] & 1'b1;
			partial_clause[0][144] 	= partial_clause_prev[0][144] & x[39];
			partial_clause[0][145] 	= partial_clause_prev[0][145] & 1'b1;
			partial_clause[0][146] 	= partial_clause_prev[0][146] & 1'b1;
			partial_clause[0][147] 	= partial_clause_prev[0][147] & 1'b1;
			partial_clause[0][148] 	= partial_clause_prev[0][148] & 1'b1;
			partial_clause[0][149] 	= partial_clause_prev[0][149] & 1'b1;
			partial_clause[0][150] 	= partial_clause_prev[0][150] & 1'b1;
			partial_clause[0][151] 	= partial_clause_prev[0][151] & 1'b1;
			partial_clause[0][152] 	= partial_clause_prev[0][152] & 1'b1;
			partial_clause[0][153] 	= partial_clause_prev[0][153] & 1'b1;
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & 1'b1;
			partial_clause[0][156] 	= partial_clause_prev[0][156] & 1'b1;
			partial_clause[0][157] 	= partial_clause_prev[0][157] & 1'b1;
			partial_clause[0][158] 	= partial_clause_prev[0][158] & 1'b1;
			partial_clause[0][159] 	= partial_clause_prev[0][159] & 1'b1;
			partial_clause[0][160] 	= partial_clause_prev[0][160] & 1'b1;
			partial_clause[0][161] 	= partial_clause_prev[0][161] & 1'b1;
			partial_clause[0][162] 	= partial_clause_prev[0][162] & 1'b1;
			partial_clause[0][163] 	= partial_clause_prev[0][163] & 1'b1;
			partial_clause[0][164] 	= partial_clause_prev[0][164] & 1'b1;
			partial_clause[0][165] 	= partial_clause_prev[0][165] & 1'b1;
			partial_clause[0][166] 	= partial_clause_prev[0][166] & 1'b1;
			partial_clause[0][167] 	= partial_clause_prev[0][167] & 1'b1;
			partial_clause[0][168] 	= partial_clause_prev[0][168] & 1'b1;
			partial_clause[0][169] 	= partial_clause_prev[0][169] & 1'b1;
			partial_clause[0][170] 	= partial_clause_prev[0][170] & 1'b1;
			partial_clause[0][171] 	= partial_clause_prev[0][171] & 1'b1;
			partial_clause[0][172] 	= partial_clause_prev[0][172] & 1'b1;
			partial_clause[0][173] 	= partial_clause_prev[0][173] & 1'b1;
			partial_clause[0][174] 	= partial_clause_prev[0][174] & 1'b1;
			partial_clause[0][175] 	= partial_clause_prev[0][175] & 1'b1;
			partial_clause[0][176] 	= partial_clause_prev[0][176] & 1'b1;
			partial_clause[0][177] 	= partial_clause_prev[0][177] & 1'b1;
			partial_clause[0][178] 	= partial_clause_prev[0][178] & x[57];
			partial_clause[0][179] 	= partial_clause_prev[0][179] & 1'b1;
			partial_clause[0][180] 	= partial_clause_prev[0][180] & 1'b1;
			partial_clause[0][181] 	= partial_clause_prev[0][181] & 1'b1;
			partial_clause[0][182] 	= partial_clause_prev[0][182] & 1'b1;
			partial_clause[0][183] 	= partial_clause_prev[0][183] & 1'b1;
			partial_clause[0][184] 	= partial_clause_prev[0][184] & 1'b1;
			partial_clause[0][185] 	= partial_clause_prev[0][185] & 1'b1;
			partial_clause[0][186] 	= partial_clause_prev[0][186] & 1'b1;
			partial_clause[0][187] 	= partial_clause_prev[0][187] & 1'b1;
			partial_clause[0][188] 	= partial_clause_prev[0][188] & 1'b1;
			partial_clause[0][189] 	= partial_clause_prev[0][189] & 1'b1;
			partial_clause[0][190] 	= partial_clause_prev[0][190] & 1'b1;
			partial_clause[0][191] 	= partial_clause_prev[0][191] & 1'b1;
			partial_clause[0][192] 	= partial_clause_prev[0][192] & 1'b1;
			partial_clause[0][193] 	= partial_clause_prev[0][193] & 1'b1;
			partial_clause[0][194] 	= partial_clause_prev[0][194] & 1'b1;
			partial_clause[0][195] 	= partial_clause_prev[0][195] & 1'b1;
			partial_clause[0][196] 	= partial_clause_prev[0][196] & 1'b1;
			partial_clause[0][197] 	= partial_clause_prev[0][197] & 1'b1;
			partial_clause[0][198] 	= partial_clause_prev[0][198] & 1'b1;
			partial_clause[0][199] 	= partial_clause_prev[0][199] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & x[56];
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & x[53];
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & x[27];
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & x[47];
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & x[4];
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & ~x[62];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & x[43];
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & x[48];
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & 1'b1;
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & ~x[62];
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			partial_clause[1][100] 	= partial_clause_prev[1][100] & 1'b1;
			partial_clause[1][101] 	= partial_clause_prev[1][101] & 1'b1;
			partial_clause[1][102] 	= partial_clause_prev[1][102] & 1'b1;
			partial_clause[1][103] 	= partial_clause_prev[1][103] & 1'b1;
			partial_clause[1][104] 	= partial_clause_prev[1][104] & 1'b1;
			partial_clause[1][105] 	= partial_clause_prev[1][105] & 1'b1;
			partial_clause[1][106] 	= partial_clause_prev[1][106] & 1'b1;
			partial_clause[1][107] 	= partial_clause_prev[1][107] & 1'b1;
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & 1'b1;
			partial_clause[1][110] 	= partial_clause_prev[1][110] & 1'b1;
			partial_clause[1][111] 	= partial_clause_prev[1][111] & 1'b1;
			partial_clause[1][112] 	= partial_clause_prev[1][112] & 1'b1;
			partial_clause[1][113] 	= partial_clause_prev[1][113] & 1'b1;
			partial_clause[1][114] 	= partial_clause_prev[1][114] & 1'b1;
			partial_clause[1][115] 	= partial_clause_prev[1][115] & 1'b1;
			partial_clause[1][116] 	= partial_clause_prev[1][116] & 1'b1;
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & 1'b1;
			partial_clause[1][119] 	= partial_clause_prev[1][119] & 1'b1;
			partial_clause[1][120] 	= partial_clause_prev[1][120] & ~x[60] & ~x[61];
			partial_clause[1][121] 	= partial_clause_prev[1][121] & 1'b1;
			partial_clause[1][122] 	= partial_clause_prev[1][122] & 1'b1;
			partial_clause[1][123] 	= partial_clause_prev[1][123] & 1'b1;
			partial_clause[1][124] 	= partial_clause_prev[1][124] & 1'b1;
			partial_clause[1][125] 	= partial_clause_prev[1][125] & ~x[63];
			partial_clause[1][126] 	= partial_clause_prev[1][126] & 1'b1;
			partial_clause[1][127] 	= partial_clause_prev[1][127] & 1'b1;
			partial_clause[1][128] 	= partial_clause_prev[1][128] & 1'b1;
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & 1'b1;
			partial_clause[1][131] 	= partial_clause_prev[1][131] & 1'b1;
			partial_clause[1][132] 	= partial_clause_prev[1][132] & 1'b1;
			partial_clause[1][133] 	= partial_clause_prev[1][133] & 1'b1;
			partial_clause[1][134] 	= partial_clause_prev[1][134] & 1'b1;
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & 1'b1;
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & 1'b1;
			partial_clause[1][139] 	= partial_clause_prev[1][139] & 1'b1;
			partial_clause[1][140] 	= partial_clause_prev[1][140] & 1'b1;
			partial_clause[1][141] 	= partial_clause_prev[1][141] & 1'b1;
			partial_clause[1][142] 	= partial_clause_prev[1][142] & 1'b1;
			partial_clause[1][143] 	= partial_clause_prev[1][143] & 1'b1;
			partial_clause[1][144] 	= partial_clause_prev[1][144] & 1'b1;
			partial_clause[1][145] 	= partial_clause_prev[1][145] & 1'b1;
			partial_clause[1][146] 	= partial_clause_prev[1][146] & 1'b1;
			partial_clause[1][147] 	= partial_clause_prev[1][147] & ~x[36] & ~x[37];
			partial_clause[1][148] 	= partial_clause_prev[1][148] & 1'b1;
			partial_clause[1][149] 	= partial_clause_prev[1][149] & 1'b1;
			partial_clause[1][150] 	= partial_clause_prev[1][150] & ~x[15];
			partial_clause[1][151] 	= partial_clause_prev[1][151] & 1'b1;
			partial_clause[1][152] 	= partial_clause_prev[1][152] & 1'b1;
			partial_clause[1][153] 	= partial_clause_prev[1][153] & 1'b1;
			partial_clause[1][154] 	= partial_clause_prev[1][154] & 1'b1;
			partial_clause[1][155] 	= partial_clause_prev[1][155] & 1'b1;
			partial_clause[1][156] 	= partial_clause_prev[1][156] & 1'b1;
			partial_clause[1][157] 	= partial_clause_prev[1][157] & 1'b1;
			partial_clause[1][158] 	= partial_clause_prev[1][158] & 1'b1;
			partial_clause[1][159] 	= partial_clause_prev[1][159] & 1'b1;
			partial_clause[1][160] 	= partial_clause_prev[1][160] & ~x[63];
			partial_clause[1][161] 	= partial_clause_prev[1][161] & 1'b1;
			partial_clause[1][162] 	= partial_clause_prev[1][162] & 1'b1;
			partial_clause[1][163] 	= partial_clause_prev[1][163] & 1'b1;
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & 1'b1;
			partial_clause[1][166] 	= partial_clause_prev[1][166] & 1'b1;
			partial_clause[1][167] 	= partial_clause_prev[1][167] & 1'b1;
			partial_clause[1][168] 	= partial_clause_prev[1][168] & 1'b1;
			partial_clause[1][169] 	= partial_clause_prev[1][169] & 1'b1;
			partial_clause[1][170] 	= partial_clause_prev[1][170] & 1'b1;
			partial_clause[1][171] 	= partial_clause_prev[1][171] & 1'b1;
			partial_clause[1][172] 	= partial_clause_prev[1][172] & ~x[63];
			partial_clause[1][173] 	= partial_clause_prev[1][173] & 1'b1;
			partial_clause[1][174] 	= partial_clause_prev[1][174] & 1'b1;
			partial_clause[1][175] 	= partial_clause_prev[1][175] & 1'b1;
			partial_clause[1][176] 	= partial_clause_prev[1][176] & 1'b1;
			partial_clause[1][177] 	= partial_clause_prev[1][177] & 1'b1;
			partial_clause[1][178] 	= partial_clause_prev[1][178] & 1'b1;
			partial_clause[1][179] 	= partial_clause_prev[1][179] & 1'b1;
			partial_clause[1][180] 	= partial_clause_prev[1][180] & 1'b1;
			partial_clause[1][181] 	= partial_clause_prev[1][181] & 1'b1;
			partial_clause[1][182] 	= partial_clause_prev[1][182] & 1'b1;
			partial_clause[1][183] 	= partial_clause_prev[1][183] & 1'b1;
			partial_clause[1][184] 	= partial_clause_prev[1][184] & 1'b1;
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & 1'b1;
			partial_clause[1][187] 	= partial_clause_prev[1][187] & 1'b1;
			partial_clause[1][188] 	= partial_clause_prev[1][188] & 1'b1;
			partial_clause[1][189] 	= partial_clause_prev[1][189] & 1'b1;
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & 1'b1;
			partial_clause[1][192] 	= partial_clause_prev[1][192] & 1'b1;
			partial_clause[1][193] 	= partial_clause_prev[1][193] & 1'b1;
			partial_clause[1][194] 	= partial_clause_prev[1][194] & 1'b1;
			partial_clause[1][195] 	= partial_clause_prev[1][195] & 1'b1;
			partial_clause[1][196] 	= partial_clause_prev[1][196] & 1'b1;
			partial_clause[1][197] 	= partial_clause_prev[1][197] & 1'b1;
			partial_clause[1][198] 	= partial_clause_prev[1][198] & 1'b1;
			partial_clause[1][199] 	= partial_clause_prev[1][199] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & x[60];
			partial_clause[2][24] 	= partial_clause_prev[2][24] & x[63];
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & x[59];
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & x[61];
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & x[0];
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & 1'b1;
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & x[61];
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & x[31];
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			partial_clause[2][100] 	= partial_clause_prev[2][100] & 1'b1;
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & 1'b1;
			partial_clause[2][103] 	= partial_clause_prev[2][103] & 1'b1;
			partial_clause[2][104] 	= partial_clause_prev[2][104] & 1'b1;
			partial_clause[2][105] 	= partial_clause_prev[2][105] & 1'b1;
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & 1'b1;
			partial_clause[2][108] 	= partial_clause_prev[2][108] & 1'b1;
			partial_clause[2][109] 	= partial_clause_prev[2][109] & 1'b1;
			partial_clause[2][110] 	= partial_clause_prev[2][110] & 1'b1;
			partial_clause[2][111] 	= partial_clause_prev[2][111] & 1'b1;
			partial_clause[2][112] 	= partial_clause_prev[2][112] & 1'b1;
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & 1'b1;
			partial_clause[2][115] 	= partial_clause_prev[2][115] & 1'b1;
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & 1'b1;
			partial_clause[2][118] 	= partial_clause_prev[2][118] & 1'b1;
			partial_clause[2][119] 	= partial_clause_prev[2][119] & 1'b1;
			partial_clause[2][120] 	= partial_clause_prev[2][120] & 1'b1;
			partial_clause[2][121] 	= partial_clause_prev[2][121] & ~x[35];
			partial_clause[2][122] 	= partial_clause_prev[2][122] & 1'b1;
			partial_clause[2][123] 	= partial_clause_prev[2][123] & 1'b1;
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & 1'b1;
			partial_clause[2][126] 	= partial_clause_prev[2][126] & 1'b1;
			partial_clause[2][127] 	= partial_clause_prev[2][127] & 1'b1;
			partial_clause[2][128] 	= partial_clause_prev[2][128] & 1'b1;
			partial_clause[2][129] 	= partial_clause_prev[2][129] & 1'b1;
			partial_clause[2][130] 	= partial_clause_prev[2][130] & 1'b1;
			partial_clause[2][131] 	= partial_clause_prev[2][131] & 1'b1;
			partial_clause[2][132] 	= partial_clause_prev[2][132] & 1'b1;
			partial_clause[2][133] 	= partial_clause_prev[2][133] & 1'b1;
			partial_clause[2][134] 	= partial_clause_prev[2][134] & 1'b1;
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & 1'b1;
			partial_clause[2][137] 	= partial_clause_prev[2][137] & 1'b1;
			partial_clause[2][138] 	= partial_clause_prev[2][138] & x[6];
			partial_clause[2][139] 	= partial_clause_prev[2][139] & x[40];
			partial_clause[2][140] 	= partial_clause_prev[2][140] & 1'b1;
			partial_clause[2][141] 	= partial_clause_prev[2][141] & 1'b1;
			partial_clause[2][142] 	= partial_clause_prev[2][142] & 1'b1;
			partial_clause[2][143] 	= partial_clause_prev[2][143] & 1'b1;
			partial_clause[2][144] 	= partial_clause_prev[2][144] & 1'b1;
			partial_clause[2][145] 	= partial_clause_prev[2][145] & 1'b1;
			partial_clause[2][146] 	= partial_clause_prev[2][146] & 1'b1;
			partial_clause[2][147] 	= partial_clause_prev[2][147] & 1'b1;
			partial_clause[2][148] 	= partial_clause_prev[2][148] & ~x[35];
			partial_clause[2][149] 	= partial_clause_prev[2][149] & 1'b1;
			partial_clause[2][150] 	= partial_clause_prev[2][150] & 1'b1;
			partial_clause[2][151] 	= partial_clause_prev[2][151] & 1'b1;
			partial_clause[2][152] 	= partial_clause_prev[2][152] & 1'b1;
			partial_clause[2][153] 	= partial_clause_prev[2][153] & 1'b1;
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & 1'b1;
			partial_clause[2][156] 	= partial_clause_prev[2][156] & 1'b1;
			partial_clause[2][157] 	= partial_clause_prev[2][157] & 1'b1;
			partial_clause[2][158] 	= partial_clause_prev[2][158] & 1'b1;
			partial_clause[2][159] 	= partial_clause_prev[2][159] & 1'b1;
			partial_clause[2][160] 	= partial_clause_prev[2][160] & 1'b1;
			partial_clause[2][161] 	= partial_clause_prev[2][161] & 1'b1;
			partial_clause[2][162] 	= partial_clause_prev[2][162] & 1'b1;
			partial_clause[2][163] 	= partial_clause_prev[2][163] & 1'b1;
			partial_clause[2][164] 	= partial_clause_prev[2][164] & 1'b1;
			partial_clause[2][165] 	= partial_clause_prev[2][165] & 1'b1;
			partial_clause[2][166] 	= partial_clause_prev[2][166] & 1'b1;
			partial_clause[2][167] 	= partial_clause_prev[2][167] & 1'b1;
			partial_clause[2][168] 	= partial_clause_prev[2][168] & 1'b1;
			partial_clause[2][169] 	= partial_clause_prev[2][169] & 1'b1;
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & 1'b1;
			partial_clause[2][173] 	= partial_clause_prev[2][173] & 1'b1;
			partial_clause[2][174] 	= partial_clause_prev[2][174] & 1'b1;
			partial_clause[2][175] 	= partial_clause_prev[2][175] & 1'b1;
			partial_clause[2][176] 	= partial_clause_prev[2][176] & 1'b1;
			partial_clause[2][177] 	= partial_clause_prev[2][177] & 1'b1;
			partial_clause[2][178] 	= partial_clause_prev[2][178] & 1'b1;
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & 1'b1;
			partial_clause[2][181] 	= partial_clause_prev[2][181] & 1'b1;
			partial_clause[2][182] 	= partial_clause_prev[2][182] & 1'b1;
			partial_clause[2][183] 	= partial_clause_prev[2][183] & 1'b1;
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & 1'b1;
			partial_clause[2][186] 	= partial_clause_prev[2][186] & 1'b1;
			partial_clause[2][187] 	= partial_clause_prev[2][187] & 1'b1;
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & 1'b1;
			partial_clause[2][190] 	= partial_clause_prev[2][190] & 1'b1;
			partial_clause[2][191] 	= partial_clause_prev[2][191] & 1'b1;
			partial_clause[2][192] 	= partial_clause_prev[2][192] & 1'b1;
			partial_clause[2][193] 	= partial_clause_prev[2][193] & 1'b1;
			partial_clause[2][194] 	= partial_clause_prev[2][194] & 1'b1;
			partial_clause[2][195] 	= partial_clause_prev[2][195] & 1'b1;
			partial_clause[2][196] 	= partial_clause_prev[2][196] & 1'b1;
			partial_clause[2][197] 	= partial_clause_prev[2][197] & 1'b1;
			partial_clause[2][198] 	= partial_clause_prev[2][198] & 1'b1;
			partial_clause[2][199] 	= partial_clause_prev[2][199] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & x[54];
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & x[48];
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & 1'b1;
			partial_clause[3][66] 	= partial_clause_prev[3][66] & x[28];
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			partial_clause[3][100] 	= partial_clause_prev[3][100] & 1'b1;
			partial_clause[3][101] 	= partial_clause_prev[3][101] & 1'b1;
			partial_clause[3][102] 	= partial_clause_prev[3][102] & 1'b1;
			partial_clause[3][103] 	= partial_clause_prev[3][103] & 1'b1;
			partial_clause[3][104] 	= partial_clause_prev[3][104] & 1'b1;
			partial_clause[3][105] 	= partial_clause_prev[3][105] & 1'b1;
			partial_clause[3][106] 	= partial_clause_prev[3][106] & 1'b1;
			partial_clause[3][107] 	= partial_clause_prev[3][107] & 1'b1;
			partial_clause[3][108] 	= partial_clause_prev[3][108] & 1'b1;
			partial_clause[3][109] 	= partial_clause_prev[3][109] & 1'b1;
			partial_clause[3][110] 	= partial_clause_prev[3][110] & 1'b1;
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & 1'b1;
			partial_clause[3][113] 	= partial_clause_prev[3][113] & 1'b1;
			partial_clause[3][114] 	= partial_clause_prev[3][114] & 1'b1;
			partial_clause[3][115] 	= partial_clause_prev[3][115] & 1'b1;
			partial_clause[3][116] 	= partial_clause_prev[3][116] & 1'b1;
			partial_clause[3][117] 	= partial_clause_prev[3][117] & 1'b1;
			partial_clause[3][118] 	= partial_clause_prev[3][118] & 1'b1;
			partial_clause[3][119] 	= partial_clause_prev[3][119] & 1'b1;
			partial_clause[3][120] 	= partial_clause_prev[3][120] & 1'b1;
			partial_clause[3][121] 	= partial_clause_prev[3][121] & 1'b1;
			partial_clause[3][122] 	= partial_clause_prev[3][122] & 1'b1;
			partial_clause[3][123] 	= partial_clause_prev[3][123] & 1'b1;
			partial_clause[3][124] 	= partial_clause_prev[3][124] & 1'b1;
			partial_clause[3][125] 	= partial_clause_prev[3][125] & 1'b1;
			partial_clause[3][126] 	= partial_clause_prev[3][126] & 1'b1;
			partial_clause[3][127] 	= partial_clause_prev[3][127] & 1'b1;
			partial_clause[3][128] 	= partial_clause_prev[3][128] & ~x[58];
			partial_clause[3][129] 	= partial_clause_prev[3][129] & 1'b1;
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & 1'b1;
			partial_clause[3][132] 	= partial_clause_prev[3][132] & 1'b1;
			partial_clause[3][133] 	= partial_clause_prev[3][133] & 1'b1;
			partial_clause[3][134] 	= partial_clause_prev[3][134] & x[13];
			partial_clause[3][135] 	= partial_clause_prev[3][135] & 1'b1;
			partial_clause[3][136] 	= partial_clause_prev[3][136] & 1'b1;
			partial_clause[3][137] 	= partial_clause_prev[3][137] & 1'b1;
			partial_clause[3][138] 	= partial_clause_prev[3][138] & 1'b1;
			partial_clause[3][139] 	= partial_clause_prev[3][139] & 1'b1;
			partial_clause[3][140] 	= partial_clause_prev[3][140] & 1'b1;
			partial_clause[3][141] 	= partial_clause_prev[3][141] & 1'b1;
			partial_clause[3][142] 	= partial_clause_prev[3][142] & 1'b1;
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & 1'b1;
			partial_clause[3][145] 	= partial_clause_prev[3][145] & 1'b1;
			partial_clause[3][146] 	= partial_clause_prev[3][146] & 1'b1;
			partial_clause[3][147] 	= partial_clause_prev[3][147] & ~x[33];
			partial_clause[3][148] 	= partial_clause_prev[3][148] & 1'b1;
			partial_clause[3][149] 	= partial_clause_prev[3][149] & 1'b1;
			partial_clause[3][150] 	= partial_clause_prev[3][150] & 1'b1;
			partial_clause[3][151] 	= partial_clause_prev[3][151] & 1'b1;
			partial_clause[3][152] 	= partial_clause_prev[3][152] & 1'b1;
			partial_clause[3][153] 	= partial_clause_prev[3][153] & 1'b1;
			partial_clause[3][154] 	= partial_clause_prev[3][154] & 1'b1;
			partial_clause[3][155] 	= partial_clause_prev[3][155] & 1'b1;
			partial_clause[3][156] 	= partial_clause_prev[3][156] & 1'b1;
			partial_clause[3][157] 	= partial_clause_prev[3][157] & 1'b1;
			partial_clause[3][158] 	= partial_clause_prev[3][158] & 1'b1;
			partial_clause[3][159] 	= partial_clause_prev[3][159] & 1'b1;
			partial_clause[3][160] 	= partial_clause_prev[3][160] & 1'b1;
			partial_clause[3][161] 	= partial_clause_prev[3][161] & 1'b1;
			partial_clause[3][162] 	= partial_clause_prev[3][162] & 1'b1;
			partial_clause[3][163] 	= partial_clause_prev[3][163] & 1'b1;
			partial_clause[3][164] 	= partial_clause_prev[3][164] & 1'b1;
			partial_clause[3][165] 	= partial_clause_prev[3][165] & 1'b1;
			partial_clause[3][166] 	= partial_clause_prev[3][166] & 1'b1;
			partial_clause[3][167] 	= partial_clause_prev[3][167] & 1'b1;
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & 1'b1;
			partial_clause[3][170] 	= partial_clause_prev[3][170] & 1'b1;
			partial_clause[3][171] 	= partial_clause_prev[3][171] & 1'b1;
			partial_clause[3][172] 	= partial_clause_prev[3][172] & 1'b1;
			partial_clause[3][173] 	= partial_clause_prev[3][173] & 1'b1;
			partial_clause[3][174] 	= partial_clause_prev[3][174] & 1'b1;
			partial_clause[3][175] 	= partial_clause_prev[3][175] & 1'b1;
			partial_clause[3][176] 	= partial_clause_prev[3][176] & 1'b1;
			partial_clause[3][177] 	= partial_clause_prev[3][177] & ~x[58];
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & 1'b1;
			partial_clause[3][180] 	= partial_clause_prev[3][180] & 1'b1;
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & 1'b1;
			partial_clause[3][183] 	= partial_clause_prev[3][183] & 1'b1;
			partial_clause[3][184] 	= partial_clause_prev[3][184] & 1'b1;
			partial_clause[3][185] 	= partial_clause_prev[3][185] & 1'b1;
			partial_clause[3][186] 	= partial_clause_prev[3][186] & ~x[60] & ~x[63];
			partial_clause[3][187] 	= partial_clause_prev[3][187] & 1'b1;
			partial_clause[3][188] 	= partial_clause_prev[3][188] & 1'b1;
			partial_clause[3][189] 	= partial_clause_prev[3][189] & 1'b1;
			partial_clause[3][190] 	= partial_clause_prev[3][190] & 1'b1;
			partial_clause[3][191] 	= partial_clause_prev[3][191] & 1'b1;
			partial_clause[3][192] 	= partial_clause_prev[3][192] & 1'b1;
			partial_clause[3][193] 	= partial_clause_prev[3][193] & 1'b1;
			partial_clause[3][194] 	= partial_clause_prev[3][194] & ~x[59] & ~x[62];
			partial_clause[3][195] 	= partial_clause_prev[3][195] & 1'b1;
			partial_clause[3][196] 	= partial_clause_prev[3][196] & 1'b1;
			partial_clause[3][197] 	= partial_clause_prev[3][197] & 1'b1;
			partial_clause[3][198] 	= partial_clause_prev[3][198] & 1'b1;
			partial_clause[3][199] 	= partial_clause_prev[3][199] & ~x[60];
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & ~x[34];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & x[45];
			partial_clause[4][12] 	= partial_clause_prev[4][12] & x[23];
			partial_clause[4][13] 	= partial_clause_prev[4][13] & ~x[32] & ~x[33];
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & ~x[34];
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & x[52];
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & x[16];
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & ~x[33];
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & x[44];
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & x[53];
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[63];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[62];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & ~x[31] & ~x[35];
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & ~x[30] & ~x[34];
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & x[55];
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & ~x[31];
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & ~x[32];
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & ~x[57] & ~x[63];
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & ~x[61];
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & ~x[58];
			partial_clause[4][91] 	= partial_clause_prev[4][91] & ~x[34];
			partial_clause[4][92] 	= partial_clause_prev[4][92] & x[46];
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & ~x[62];
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			partial_clause[4][100] 	= partial_clause_prev[4][100] & x[32];
			partial_clause[4][101] 	= partial_clause_prev[4][101] & x[37];
			partial_clause[4][102] 	= partial_clause_prev[4][102] & 1'b1;
			partial_clause[4][103] 	= partial_clause_prev[4][103] & 1'b1;
			partial_clause[4][104] 	= partial_clause_prev[4][104] & 1'b1;
			partial_clause[4][105] 	= partial_clause_prev[4][105] & 1'b1;
			partial_clause[4][106] 	= partial_clause_prev[4][106] & 1'b1;
			partial_clause[4][107] 	= partial_clause_prev[4][107] & 1'b1;
			partial_clause[4][108] 	= partial_clause_prev[4][108] & 1'b1;
			partial_clause[4][109] 	= partial_clause_prev[4][109] & 1'b1;
			partial_clause[4][110] 	= partial_clause_prev[4][110] & 1'b1;
			partial_clause[4][111] 	= partial_clause_prev[4][111] & 1'b1;
			partial_clause[4][112] 	= partial_clause_prev[4][112] & x[61];
			partial_clause[4][113] 	= partial_clause_prev[4][113] & 1'b1;
			partial_clause[4][114] 	= partial_clause_prev[4][114] & 1'b1;
			partial_clause[4][115] 	= partial_clause_prev[4][115] & x[31];
			partial_clause[4][116] 	= partial_clause_prev[4][116] & 1'b1;
			partial_clause[4][117] 	= partial_clause_prev[4][117] & ~x[26];
			partial_clause[4][118] 	= partial_clause_prev[4][118] & 1'b1;
			partial_clause[4][119] 	= partial_clause_prev[4][119] & 1'b1;
			partial_clause[4][120] 	= partial_clause_prev[4][120] & 1'b1;
			partial_clause[4][121] 	= partial_clause_prev[4][121] & 1'b1;
			partial_clause[4][122] 	= partial_clause_prev[4][122] & 1'b1;
			partial_clause[4][123] 	= partial_clause_prev[4][123] & x[38];
			partial_clause[4][124] 	= partial_clause_prev[4][124] & 1'b1;
			partial_clause[4][125] 	= partial_clause_prev[4][125] & 1'b1;
			partial_clause[4][126] 	= partial_clause_prev[4][126] & 1'b1;
			partial_clause[4][127] 	= partial_clause_prev[4][127] & 1'b1;
			partial_clause[4][128] 	= partial_clause_prev[4][128] & 1'b1;
			partial_clause[4][129] 	= partial_clause_prev[4][129] & 1'b1;
			partial_clause[4][130] 	= partial_clause_prev[4][130] & 1'b1;
			partial_clause[4][131] 	= partial_clause_prev[4][131] & 1'b1;
			partial_clause[4][132] 	= partial_clause_prev[4][132] & 1'b1;
			partial_clause[4][133] 	= partial_clause_prev[4][133] & 1'b1;
			partial_clause[4][134] 	= partial_clause_prev[4][134] & 1'b1;
			partial_clause[4][135] 	= partial_clause_prev[4][135] & 1'b1;
			partial_clause[4][136] 	= partial_clause_prev[4][136] & 1'b1;
			partial_clause[4][137] 	= partial_clause_prev[4][137] & 1'b1;
			partial_clause[4][138] 	= partial_clause_prev[4][138] & 1'b1;
			partial_clause[4][139] 	= partial_clause_prev[4][139] & 1'b1;
			partial_clause[4][140] 	= partial_clause_prev[4][140] & 1'b1;
			partial_clause[4][141] 	= partial_clause_prev[4][141] & 1'b1;
			partial_clause[4][142] 	= partial_clause_prev[4][142] & 1'b1;
			partial_clause[4][143] 	= partial_clause_prev[4][143] & 1'b1;
			partial_clause[4][144] 	= partial_clause_prev[4][144] & 1'b1;
			partial_clause[4][145] 	= partial_clause_prev[4][145] & 1'b1;
			partial_clause[4][146] 	= partial_clause_prev[4][146] & 1'b1;
			partial_clause[4][147] 	= partial_clause_prev[4][147] & 1'b1;
			partial_clause[4][148] 	= partial_clause_prev[4][148] & 1'b1;
			partial_clause[4][149] 	= partial_clause_prev[4][149] & x[63];
			partial_clause[4][150] 	= partial_clause_prev[4][150] & 1'b1;
			partial_clause[4][151] 	= partial_clause_prev[4][151] & 1'b1;
			partial_clause[4][152] 	= partial_clause_prev[4][152] & 1'b1;
			partial_clause[4][153] 	= partial_clause_prev[4][153] & 1'b1;
			partial_clause[4][154] 	= partial_clause_prev[4][154] & 1'b1;
			partial_clause[4][155] 	= partial_clause_prev[4][155] & 1'b1;
			partial_clause[4][156] 	= partial_clause_prev[4][156] & 1'b1;
			partial_clause[4][157] 	= partial_clause_prev[4][157] & 1'b1;
			partial_clause[4][158] 	= partial_clause_prev[4][158] & 1'b1;
			partial_clause[4][159] 	= partial_clause_prev[4][159] & 1'b1;
			partial_clause[4][160] 	= partial_clause_prev[4][160] & 1'b1;
			partial_clause[4][161] 	= partial_clause_prev[4][161] & ~x[11];
			partial_clause[4][162] 	= partial_clause_prev[4][162] & 1'b1;
			partial_clause[4][163] 	= partial_clause_prev[4][163] & 1'b1;
			partial_clause[4][164] 	= partial_clause_prev[4][164] & 1'b1;
			partial_clause[4][165] 	= partial_clause_prev[4][165] & 1'b1;
			partial_clause[4][166] 	= partial_clause_prev[4][166] & 1'b1;
			partial_clause[4][167] 	= partial_clause_prev[4][167] & 1'b1;
			partial_clause[4][168] 	= partial_clause_prev[4][168] & 1'b1;
			partial_clause[4][169] 	= partial_clause_prev[4][169] & 1'b1;
			partial_clause[4][170] 	= partial_clause_prev[4][170] & 1'b1;
			partial_clause[4][171] 	= partial_clause_prev[4][171] & 1'b1;
			partial_clause[4][172] 	= partial_clause_prev[4][172] & 1'b1;
			partial_clause[4][173] 	= partial_clause_prev[4][173] & x[36];
			partial_clause[4][174] 	= partial_clause_prev[4][174] & 1'b1;
			partial_clause[4][175] 	= partial_clause_prev[4][175] & x[60];
			partial_clause[4][176] 	= partial_clause_prev[4][176] & 1'b1;
			partial_clause[4][177] 	= partial_clause_prev[4][177] & 1'b1;
			partial_clause[4][178] 	= partial_clause_prev[4][178] & 1'b1;
			partial_clause[4][179] 	= partial_clause_prev[4][179] & x[60];
			partial_clause[4][180] 	= partial_clause_prev[4][180] & 1'b1;
			partial_clause[4][181] 	= partial_clause_prev[4][181] & 1'b1;
			partial_clause[4][182] 	= partial_clause_prev[4][182] & 1'b1;
			partial_clause[4][183] 	= partial_clause_prev[4][183] & 1'b1;
			partial_clause[4][184] 	= partial_clause_prev[4][184] & 1'b1;
			partial_clause[4][185] 	= partial_clause_prev[4][185] & 1'b1;
			partial_clause[4][186] 	= partial_clause_prev[4][186] & 1'b1;
			partial_clause[4][187] 	= partial_clause_prev[4][187] & 1'b1;
			partial_clause[4][188] 	= partial_clause_prev[4][188] & 1'b1;
			partial_clause[4][189] 	= partial_clause_prev[4][189] & 1'b1;
			partial_clause[4][190] 	= partial_clause_prev[4][190] & 1'b1;
			partial_clause[4][191] 	= partial_clause_prev[4][191] & 1'b1;
			partial_clause[4][192] 	= partial_clause_prev[4][192] & 1'b1;
			partial_clause[4][193] 	= partial_clause_prev[4][193] & 1'b1;
			partial_clause[4][194] 	= partial_clause_prev[4][194] & 1'b1;
			partial_clause[4][195] 	= partial_clause_prev[4][195] & 1'b1;
			partial_clause[4][196] 	= partial_clause_prev[4][196] & 1'b1;
			partial_clause[4][197] 	= partial_clause_prev[4][197] & 1'b1;
			partial_clause[4][198] 	= partial_clause_prev[4][198] & 1'b1;
			partial_clause[4][199] 	= partial_clause_prev[4][199] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & ~x[7];
			partial_clause[5][12] 	= partial_clause_prev[5][12] & ~x[36];
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & x[25];
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & ~x[60];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & ~x[34];
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & ~x[61];
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & x[42];
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			partial_clause[5][100] 	= partial_clause_prev[5][100] & 1'b1;
			partial_clause[5][101] 	= partial_clause_prev[5][101] & 1'b1;
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & 1'b1;
			partial_clause[5][104] 	= partial_clause_prev[5][104] & x[57];
			partial_clause[5][105] 	= partial_clause_prev[5][105] & 1'b1;
			partial_clause[5][106] 	= partial_clause_prev[5][106] & 1'b1;
			partial_clause[5][107] 	= partial_clause_prev[5][107] & 1'b1;
			partial_clause[5][108] 	= partial_clause_prev[5][108] & 1'b1;
			partial_clause[5][109] 	= partial_clause_prev[5][109] & 1'b1;
			partial_clause[5][110] 	= partial_clause_prev[5][110] & 1'b1;
			partial_clause[5][111] 	= partial_clause_prev[5][111] & x[37];
			partial_clause[5][112] 	= partial_clause_prev[5][112] & 1'b1;
			partial_clause[5][113] 	= partial_clause_prev[5][113] & x[33];
			partial_clause[5][114] 	= partial_clause_prev[5][114] & 1'b1;
			partial_clause[5][115] 	= partial_clause_prev[5][115] & 1'b1;
			partial_clause[5][116] 	= partial_clause_prev[5][116] & 1'b1;
			partial_clause[5][117] 	= partial_clause_prev[5][117] & 1'b1;
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & 1'b1;
			partial_clause[5][120] 	= partial_clause_prev[5][120] & 1'b1;
			partial_clause[5][121] 	= partial_clause_prev[5][121] & 1'b1;
			partial_clause[5][122] 	= partial_clause_prev[5][122] & 1'b1;
			partial_clause[5][123] 	= partial_clause_prev[5][123] & 1'b1;
			partial_clause[5][124] 	= partial_clause_prev[5][124] & 1'b1;
			partial_clause[5][125] 	= partial_clause_prev[5][125] & 1'b1;
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & 1'b1;
			partial_clause[5][128] 	= partial_clause_prev[5][128] & 1'b1;
			partial_clause[5][129] 	= partial_clause_prev[5][129] & 1'b1;
			partial_clause[5][130] 	= partial_clause_prev[5][130] & 1'b1;
			partial_clause[5][131] 	= partial_clause_prev[5][131] & 1'b1;
			partial_clause[5][132] 	= partial_clause_prev[5][132] & 1'b1;
			partial_clause[5][133] 	= partial_clause_prev[5][133] & 1'b1;
			partial_clause[5][134] 	= partial_clause_prev[5][134] & 1'b1;
			partial_clause[5][135] 	= partial_clause_prev[5][135] & 1'b1;
			partial_clause[5][136] 	= partial_clause_prev[5][136] & 1'b1;
			partial_clause[5][137] 	= partial_clause_prev[5][137] & x[6];
			partial_clause[5][138] 	= partial_clause_prev[5][138] & x[29];
			partial_clause[5][139] 	= partial_clause_prev[5][139] & x[6];
			partial_clause[5][140] 	= partial_clause_prev[5][140] & 1'b1;
			partial_clause[5][141] 	= partial_clause_prev[5][141] & 1'b1;
			partial_clause[5][142] 	= partial_clause_prev[5][142] & 1'b1;
			partial_clause[5][143] 	= partial_clause_prev[5][143] & 1'b1;
			partial_clause[5][144] 	= partial_clause_prev[5][144] & 1'b1;
			partial_clause[5][145] 	= partial_clause_prev[5][145] & 1'b1;
			partial_clause[5][146] 	= partial_clause_prev[5][146] & 1'b1;
			partial_clause[5][147] 	= partial_clause_prev[5][147] & 1'b1;
			partial_clause[5][148] 	= partial_clause_prev[5][148] & 1'b1;
			partial_clause[5][149] 	= partial_clause_prev[5][149] & 1'b1;
			partial_clause[5][150] 	= partial_clause_prev[5][150] & 1'b1;
			partial_clause[5][151] 	= partial_clause_prev[5][151] & 1'b1;
			partial_clause[5][152] 	= partial_clause_prev[5][152] & 1'b1;
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & 1'b1;
			partial_clause[5][155] 	= partial_clause_prev[5][155] & 1'b1;
			partial_clause[5][156] 	= partial_clause_prev[5][156] & 1'b1;
			partial_clause[5][157] 	= partial_clause_prev[5][157] & 1'b1;
			partial_clause[5][158] 	= partial_clause_prev[5][158] & 1'b1;
			partial_clause[5][159] 	= partial_clause_prev[5][159] & 1'b1;
			partial_clause[5][160] 	= partial_clause_prev[5][160] & 1'b1;
			partial_clause[5][161] 	= partial_clause_prev[5][161] & 1'b1;
			partial_clause[5][162] 	= partial_clause_prev[5][162] & 1'b1;
			partial_clause[5][163] 	= partial_clause_prev[5][163] & 1'b1;
			partial_clause[5][164] 	= partial_clause_prev[5][164] & 1'b1;
			partial_clause[5][165] 	= partial_clause_prev[5][165] & 1'b1;
			partial_clause[5][166] 	= partial_clause_prev[5][166] & 1'b1;
			partial_clause[5][167] 	= partial_clause_prev[5][167] & 1'b1;
			partial_clause[5][168] 	= partial_clause_prev[5][168] & 1'b1;
			partial_clause[5][169] 	= partial_clause_prev[5][169] & 1'b1;
			partial_clause[5][170] 	= partial_clause_prev[5][170] & 1'b1;
			partial_clause[5][171] 	= partial_clause_prev[5][171] & x[6];
			partial_clause[5][172] 	= partial_clause_prev[5][172] & 1'b1;
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & 1'b1;
			partial_clause[5][175] 	= partial_clause_prev[5][175] & 1'b1;
			partial_clause[5][176] 	= partial_clause_prev[5][176] & 1'b1;
			partial_clause[5][177] 	= partial_clause_prev[5][177] & 1'b1;
			partial_clause[5][178] 	= partial_clause_prev[5][178] & 1'b1;
			partial_clause[5][179] 	= partial_clause_prev[5][179] & 1'b1;
			partial_clause[5][180] 	= partial_clause_prev[5][180] & 1'b1;
			partial_clause[5][181] 	= partial_clause_prev[5][181] & 1'b1;
			partial_clause[5][182] 	= partial_clause_prev[5][182] & 1'b1;
			partial_clause[5][183] 	= partial_clause_prev[5][183] & 1'b1;
			partial_clause[5][184] 	= partial_clause_prev[5][184] & 1'b1;
			partial_clause[5][185] 	= partial_clause_prev[5][185] & 1'b1;
			partial_clause[5][186] 	= partial_clause_prev[5][186] & 1'b1;
			partial_clause[5][187] 	= partial_clause_prev[5][187] & ~x[38] & ~x[40];
			partial_clause[5][188] 	= partial_clause_prev[5][188] & 1'b1;
			partial_clause[5][189] 	= partial_clause_prev[5][189] & 1'b1;
			partial_clause[5][190] 	= partial_clause_prev[5][190] & 1'b1;
			partial_clause[5][191] 	= partial_clause_prev[5][191] & x[50];
			partial_clause[5][192] 	= partial_clause_prev[5][192] & 1'b1;
			partial_clause[5][193] 	= partial_clause_prev[5][193] & 1'b1;
			partial_clause[5][194] 	= partial_clause_prev[5][194] & 1'b1;
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & x[34];
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & 1'b1;
			partial_clause[5][199] 	= partial_clause_prev[5][199] & x[59];
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & ~x[62] & ~x[63];
			partial_clause[6][1] 	= partial_clause_prev[6][1] & x[20];
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & x[6];
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & ~x[63];
			partial_clause[6][23] 	= partial_clause_prev[6][23] & x[4];
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & x[44];
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & x[4];
			partial_clause[6][31] 	= partial_clause_prev[6][31] & x[41];
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & x[10];
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & x[39];
			partial_clause[6][41] 	= partial_clause_prev[6][41] & ~x[61];
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & ~x[60];
			partial_clause[6][46] 	= partial_clause_prev[6][46] & ~x[59];
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & x[10];
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & x[41];
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & x[42];
			partial_clause[6][69] 	= partial_clause_prev[6][69] & x[11];
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & x[39];
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & x[3];
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & ~x[62];
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & x[6];
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & x[5];
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & x[36];
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			partial_clause[6][100] 	= partial_clause_prev[6][100] & ~x[36] & ~x[39];
			partial_clause[6][101] 	= partial_clause_prev[6][101] & 1'b1;
			partial_clause[6][102] 	= partial_clause_prev[6][102] & 1'b1;
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & 1'b1;
			partial_clause[6][105] 	= partial_clause_prev[6][105] & 1'b1;
			partial_clause[6][106] 	= partial_clause_prev[6][106] & 1'b1;
			partial_clause[6][107] 	= partial_clause_prev[6][107] & 1'b1;
			partial_clause[6][108] 	= partial_clause_prev[6][108] & 1'b1;
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & 1'b1;
			partial_clause[6][111] 	= partial_clause_prev[6][111] & ~x[6] & ~x[36];
			partial_clause[6][112] 	= partial_clause_prev[6][112] & 1'b1;
			partial_clause[6][113] 	= partial_clause_prev[6][113] & 1'b1;
			partial_clause[6][114] 	= partial_clause_prev[6][114] & 1'b1;
			partial_clause[6][115] 	= partial_clause_prev[6][115] & 1'b1;
			partial_clause[6][116] 	= partial_clause_prev[6][116] & 1'b1;
			partial_clause[6][117] 	= partial_clause_prev[6][117] & 1'b1;
			partial_clause[6][118] 	= partial_clause_prev[6][118] & 1'b1;
			partial_clause[6][119] 	= partial_clause_prev[6][119] & 1'b1;
			partial_clause[6][120] 	= partial_clause_prev[6][120] & ~x[36] & ~x[39];
			partial_clause[6][121] 	= partial_clause_prev[6][121] & 1'b1;
			partial_clause[6][122] 	= partial_clause_prev[6][122] & 1'b1;
			partial_clause[6][123] 	= partial_clause_prev[6][123] & 1'b1;
			partial_clause[6][124] 	= partial_clause_prev[6][124] & 1'b1;
			partial_clause[6][125] 	= partial_clause_prev[6][125] & 1'b1;
			partial_clause[6][126] 	= partial_clause_prev[6][126] & 1'b1;
			partial_clause[6][127] 	= partial_clause_prev[6][127] & 1'b1;
			partial_clause[6][128] 	= partial_clause_prev[6][128] & 1'b1;
			partial_clause[6][129] 	= partial_clause_prev[6][129] & 1'b1;
			partial_clause[6][130] 	= partial_clause_prev[6][130] & 1'b1;
			partial_clause[6][131] 	= partial_clause_prev[6][131] & ~x[56];
			partial_clause[6][132] 	= partial_clause_prev[6][132] & 1'b1;
			partial_clause[6][133] 	= partial_clause_prev[6][133] & ~x[33] & ~x[37];
			partial_clause[6][134] 	= partial_clause_prev[6][134] & 1'b1;
			partial_clause[6][135] 	= partial_clause_prev[6][135] & 1'b1;
			partial_clause[6][136] 	= partial_clause_prev[6][136] & 1'b1;
			partial_clause[6][137] 	= partial_clause_prev[6][137] & ~x[56];
			partial_clause[6][138] 	= partial_clause_prev[6][138] & 1'b1;
			partial_clause[6][139] 	= partial_clause_prev[6][139] & 1'b1;
			partial_clause[6][140] 	= partial_clause_prev[6][140] & 1'b1;
			partial_clause[6][141] 	= partial_clause_prev[6][141] & 1'b1;
			partial_clause[6][142] 	= partial_clause_prev[6][142] & 1'b1;
			partial_clause[6][143] 	= partial_clause_prev[6][143] & ~x[39];
			partial_clause[6][144] 	= partial_clause_prev[6][144] & 1'b1;
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & 1'b1;
			partial_clause[6][147] 	= partial_clause_prev[6][147] & 1'b1;
			partial_clause[6][148] 	= partial_clause_prev[6][148] & 1'b1;
			partial_clause[6][149] 	= partial_clause_prev[6][149] & 1'b1;
			partial_clause[6][150] 	= partial_clause_prev[6][150] & ~x[34];
			partial_clause[6][151] 	= partial_clause_prev[6][151] & 1'b1;
			partial_clause[6][152] 	= partial_clause_prev[6][152] & 1'b1;
			partial_clause[6][153] 	= partial_clause_prev[6][153] & 1'b1;
			partial_clause[6][154] 	= partial_clause_prev[6][154] & ~x[2];
			partial_clause[6][155] 	= partial_clause_prev[6][155] & 1'b1;
			partial_clause[6][156] 	= partial_clause_prev[6][156] & 1'b1;
			partial_clause[6][157] 	= partial_clause_prev[6][157] & 1'b1;
			partial_clause[6][158] 	= partial_clause_prev[6][158] & 1'b1;
			partial_clause[6][159] 	= partial_clause_prev[6][159] & 1'b1;
			partial_clause[6][160] 	= partial_clause_prev[6][160] & 1'b1;
			partial_clause[6][161] 	= partial_clause_prev[6][161] & 1'b1;
			partial_clause[6][162] 	= partial_clause_prev[6][162] & 1'b1;
			partial_clause[6][163] 	= partial_clause_prev[6][163] & 1'b1;
			partial_clause[6][164] 	= partial_clause_prev[6][164] & 1'b1;
			partial_clause[6][165] 	= partial_clause_prev[6][165] & 1'b1;
			partial_clause[6][166] 	= partial_clause_prev[6][166] & 1'b1;
			partial_clause[6][167] 	= partial_clause_prev[6][167] & 1'b1;
			partial_clause[6][168] 	= partial_clause_prev[6][168] & ~x[35];
			partial_clause[6][169] 	= partial_clause_prev[6][169] & 1'b1;
			partial_clause[6][170] 	= partial_clause_prev[6][170] & 1'b1;
			partial_clause[6][171] 	= partial_clause_prev[6][171] & ~x[34];
			partial_clause[6][172] 	= partial_clause_prev[6][172] & 1'b1;
			partial_clause[6][173] 	= partial_clause_prev[6][173] & 1'b1;
			partial_clause[6][174] 	= partial_clause_prev[6][174] & 1'b1;
			partial_clause[6][175] 	= partial_clause_prev[6][175] & 1'b1;
			partial_clause[6][176] 	= partial_clause_prev[6][176] & 1'b1;
			partial_clause[6][177] 	= partial_clause_prev[6][177] & 1'b1;
			partial_clause[6][178] 	= partial_clause_prev[6][178] & 1'b1;
			partial_clause[6][179] 	= partial_clause_prev[6][179] & 1'b1;
			partial_clause[6][180] 	= partial_clause_prev[6][180] & 1'b1;
			partial_clause[6][181] 	= partial_clause_prev[6][181] & 1'b1;
			partial_clause[6][182] 	= partial_clause_prev[6][182] & ~x[33];
			partial_clause[6][183] 	= partial_clause_prev[6][183] & 1'b1;
			partial_clause[6][184] 	= partial_clause_prev[6][184] & 1'b1;
			partial_clause[6][185] 	= partial_clause_prev[6][185] & 1'b1;
			partial_clause[6][186] 	= partial_clause_prev[6][186] & ~x[37] & ~x[39];
			partial_clause[6][187] 	= partial_clause_prev[6][187] & ~x[29] & ~x[32] & ~x[57];
			partial_clause[6][188] 	= partial_clause_prev[6][188] & 1'b1;
			partial_clause[6][189] 	= partial_clause_prev[6][189] & 1'b1;
			partial_clause[6][190] 	= partial_clause_prev[6][190] & 1'b1;
			partial_clause[6][191] 	= partial_clause_prev[6][191] & 1'b1;
			partial_clause[6][192] 	= partial_clause_prev[6][192] & 1'b1;
			partial_clause[6][193] 	= partial_clause_prev[6][193] & 1'b1;
			partial_clause[6][194] 	= partial_clause_prev[6][194] & 1'b1;
			partial_clause[6][195] 	= partial_clause_prev[6][195] & 1'b1;
			partial_clause[6][196] 	= partial_clause_prev[6][196] & 1'b1;
			partial_clause[6][197] 	= partial_clause_prev[6][197] & 1'b1;
			partial_clause[6][198] 	= partial_clause_prev[6][198] & 1'b1;
			partial_clause[6][199] 	= partial_clause_prev[6][199] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & x[20];
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & x[21];
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & ~x[62];
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & x[40];
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			partial_clause[7][100] 	= partial_clause_prev[7][100] & 1'b1;
			partial_clause[7][101] 	= partial_clause_prev[7][101] & 1'b1;
			partial_clause[7][102] 	= partial_clause_prev[7][102] & 1'b1;
			partial_clause[7][103] 	= partial_clause_prev[7][103] & 1'b1;
			partial_clause[7][104] 	= partial_clause_prev[7][104] & 1'b1;
			partial_clause[7][105] 	= partial_clause_prev[7][105] & 1'b1;
			partial_clause[7][106] 	= partial_clause_prev[7][106] & x[63];
			partial_clause[7][107] 	= partial_clause_prev[7][107] & 1'b1;
			partial_clause[7][108] 	= partial_clause_prev[7][108] & 1'b1;
			partial_clause[7][109] 	= partial_clause_prev[7][109] & 1'b1;
			partial_clause[7][110] 	= partial_clause_prev[7][110] & 1'b1;
			partial_clause[7][111] 	= partial_clause_prev[7][111] & 1'b1;
			partial_clause[7][112] 	= partial_clause_prev[7][112] & 1'b1;
			partial_clause[7][113] 	= partial_clause_prev[7][113] & 1'b1;
			partial_clause[7][114] 	= partial_clause_prev[7][114] & 1'b1;
			partial_clause[7][115] 	= partial_clause_prev[7][115] & 1'b1;
			partial_clause[7][116] 	= partial_clause_prev[7][116] & 1'b1;
			partial_clause[7][117] 	= partial_clause_prev[7][117] & 1'b1;
			partial_clause[7][118] 	= partial_clause_prev[7][118] & 1'b1;
			partial_clause[7][119] 	= partial_clause_prev[7][119] & 1'b1;
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & 1'b1;
			partial_clause[7][123] 	= partial_clause_prev[7][123] & 1'b1;
			partial_clause[7][124] 	= partial_clause_prev[7][124] & 1'b1;
			partial_clause[7][125] 	= partial_clause_prev[7][125] & 1'b1;
			partial_clause[7][126] 	= partial_clause_prev[7][126] & 1'b1;
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & 1'b1;
			partial_clause[7][129] 	= partial_clause_prev[7][129] & 1'b1;
			partial_clause[7][130] 	= partial_clause_prev[7][130] & 1'b1;
			partial_clause[7][131] 	= partial_clause_prev[7][131] & 1'b1;
			partial_clause[7][132] 	= partial_clause_prev[7][132] & 1'b1;
			partial_clause[7][133] 	= partial_clause_prev[7][133] & 1'b1;
			partial_clause[7][134] 	= partial_clause_prev[7][134] & 1'b1;
			partial_clause[7][135] 	= partial_clause_prev[7][135] & 1'b1;
			partial_clause[7][136] 	= partial_clause_prev[7][136] & 1'b1;
			partial_clause[7][137] 	= partial_clause_prev[7][137] & 1'b1;
			partial_clause[7][138] 	= partial_clause_prev[7][138] & 1'b1;
			partial_clause[7][139] 	= partial_clause_prev[7][139] & 1'b1;
			partial_clause[7][140] 	= partial_clause_prev[7][140] & 1'b1;
			partial_clause[7][141] 	= partial_clause_prev[7][141] & 1'b1;
			partial_clause[7][142] 	= partial_clause_prev[7][142] & 1'b1;
			partial_clause[7][143] 	= partial_clause_prev[7][143] & 1'b1;
			partial_clause[7][144] 	= partial_clause_prev[7][144] & 1'b1;
			partial_clause[7][145] 	= partial_clause_prev[7][145] & 1'b1;
			partial_clause[7][146] 	= partial_clause_prev[7][146] & 1'b1;
			partial_clause[7][147] 	= partial_clause_prev[7][147] & 1'b1;
			partial_clause[7][148] 	= partial_clause_prev[7][148] & 1'b1;
			partial_clause[7][149] 	= partial_clause_prev[7][149] & 1'b1;
			partial_clause[7][150] 	= partial_clause_prev[7][150] & 1'b1;
			partial_clause[7][151] 	= partial_clause_prev[7][151] & 1'b1;
			partial_clause[7][152] 	= partial_clause_prev[7][152] & 1'b1;
			partial_clause[7][153] 	= partial_clause_prev[7][153] & 1'b1;
			partial_clause[7][154] 	= partial_clause_prev[7][154] & 1'b1;
			partial_clause[7][155] 	= partial_clause_prev[7][155] & 1'b1;
			partial_clause[7][156] 	= partial_clause_prev[7][156] & 1'b1;
			partial_clause[7][157] 	= partial_clause_prev[7][157] & 1'b1;
			partial_clause[7][158] 	= partial_clause_prev[7][158] & 1'b1;
			partial_clause[7][159] 	= partial_clause_prev[7][159] & 1'b1;
			partial_clause[7][160] 	= partial_clause_prev[7][160] & 1'b1;
			partial_clause[7][161] 	= partial_clause_prev[7][161] & 1'b1;
			partial_clause[7][162] 	= partial_clause_prev[7][162] & 1'b1;
			partial_clause[7][163] 	= partial_clause_prev[7][163] & 1'b1;
			partial_clause[7][164] 	= partial_clause_prev[7][164] & 1'b1;
			partial_clause[7][165] 	= partial_clause_prev[7][165] & 1'b1;
			partial_clause[7][166] 	= partial_clause_prev[7][166] & ~x[29];
			partial_clause[7][167] 	= partial_clause_prev[7][167] & x[58];
			partial_clause[7][168] 	= partial_clause_prev[7][168] & x[63];
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & 1'b1;
			partial_clause[7][171] 	= partial_clause_prev[7][171] & 1'b1;
			partial_clause[7][172] 	= partial_clause_prev[7][172] & 1'b1;
			partial_clause[7][173] 	= partial_clause_prev[7][173] & 1'b1;
			partial_clause[7][174] 	= partial_clause_prev[7][174] & 1'b1;
			partial_clause[7][175] 	= partial_clause_prev[7][175] & 1'b1;
			partial_clause[7][176] 	= partial_clause_prev[7][176] & 1'b1;
			partial_clause[7][177] 	= partial_clause_prev[7][177] & 1'b1;
			partial_clause[7][178] 	= partial_clause_prev[7][178] & 1'b1;
			partial_clause[7][179] 	= partial_clause_prev[7][179] & 1'b1;
			partial_clause[7][180] 	= partial_clause_prev[7][180] & 1'b1;
			partial_clause[7][181] 	= partial_clause_prev[7][181] & 1'b1;
			partial_clause[7][182] 	= partial_clause_prev[7][182] & 1'b1;
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & 1'b1;
			partial_clause[7][185] 	= partial_clause_prev[7][185] & 1'b1;
			partial_clause[7][186] 	= partial_clause_prev[7][186] & 1'b1;
			partial_clause[7][187] 	= partial_clause_prev[7][187] & 1'b1;
			partial_clause[7][188] 	= partial_clause_prev[7][188] & 1'b1;
			partial_clause[7][189] 	= partial_clause_prev[7][189] & 1'b1;
			partial_clause[7][190] 	= partial_clause_prev[7][190] & 1'b1;
			partial_clause[7][191] 	= partial_clause_prev[7][191] & 1'b1;
			partial_clause[7][192] 	= partial_clause_prev[7][192] & 1'b1;
			partial_clause[7][193] 	= partial_clause_prev[7][193] & 1'b1;
			partial_clause[7][194] 	= partial_clause_prev[7][194] & 1'b1;
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & 1'b1;
			partial_clause[7][197] 	= partial_clause_prev[7][197] & 1'b1;
			partial_clause[7][198] 	= partial_clause_prev[7][198] & 1'b1;
			partial_clause[7][199] 	= partial_clause_prev[7][199] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & ~x[35] & ~x[59];
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & x[21];
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & x[48];
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & ~x[34];
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			partial_clause[8][100] 	= partial_clause_prev[8][100] & x[35];
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & 1'b1;
			partial_clause[8][103] 	= partial_clause_prev[8][103] & 1'b1;
			partial_clause[8][104] 	= partial_clause_prev[8][104] & 1'b1;
			partial_clause[8][105] 	= partial_clause_prev[8][105] & 1'b1;
			partial_clause[8][106] 	= partial_clause_prev[8][106] & 1'b1;
			partial_clause[8][107] 	= partial_clause_prev[8][107] & 1'b1;
			partial_clause[8][108] 	= partial_clause_prev[8][108] & 1'b1;
			partial_clause[8][109] 	= partial_clause_prev[8][109] & 1'b1;
			partial_clause[8][110] 	= partial_clause_prev[8][110] & 1'b1;
			partial_clause[8][111] 	= partial_clause_prev[8][111] & 1'b1;
			partial_clause[8][112] 	= partial_clause_prev[8][112] & 1'b1;
			partial_clause[8][113] 	= partial_clause_prev[8][113] & 1'b1;
			partial_clause[8][114] 	= partial_clause_prev[8][114] & 1'b1;
			partial_clause[8][115] 	= partial_clause_prev[8][115] & 1'b1;
			partial_clause[8][116] 	= partial_clause_prev[8][116] & x[36];
			partial_clause[8][117] 	= partial_clause_prev[8][117] & 1'b1;
			partial_clause[8][118] 	= partial_clause_prev[8][118] & 1'b1;
			partial_clause[8][119] 	= partial_clause_prev[8][119] & 1'b1;
			partial_clause[8][120] 	= partial_clause_prev[8][120] & 1'b1;
			partial_clause[8][121] 	= partial_clause_prev[8][121] & x[36];
			partial_clause[8][122] 	= partial_clause_prev[8][122] & 1'b1;
			partial_clause[8][123] 	= partial_clause_prev[8][123] & 1'b1;
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & 1'b1;
			partial_clause[8][126] 	= partial_clause_prev[8][126] & 1'b1;
			partial_clause[8][127] 	= partial_clause_prev[8][127] & 1'b1;
			partial_clause[8][128] 	= partial_clause_prev[8][128] & 1'b1;
			partial_clause[8][129] 	= partial_clause_prev[8][129] & 1'b1;
			partial_clause[8][130] 	= partial_clause_prev[8][130] & 1'b1;
			partial_clause[8][131] 	= partial_clause_prev[8][131] & x[34];
			partial_clause[8][132] 	= partial_clause_prev[8][132] & ~x[60];
			partial_clause[8][133] 	= partial_clause_prev[8][133] & 1'b1;
			partial_clause[8][134] 	= partial_clause_prev[8][134] & 1'b1;
			partial_clause[8][135] 	= partial_clause_prev[8][135] & 1'b1;
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & 1'b1;
			partial_clause[8][138] 	= partial_clause_prev[8][138] & 1'b1;
			partial_clause[8][139] 	= partial_clause_prev[8][139] & 1'b1;
			partial_clause[8][140] 	= partial_clause_prev[8][140] & 1'b1;
			partial_clause[8][141] 	= partial_clause_prev[8][141] & 1'b1;
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & 1'b1;
			partial_clause[8][144] 	= partial_clause_prev[8][144] & 1'b1;
			partial_clause[8][145] 	= partial_clause_prev[8][145] & 1'b1;
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & 1'b1;
			partial_clause[8][148] 	= partial_clause_prev[8][148] & 1'b1;
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & x[5];
			partial_clause[8][151] 	= partial_clause_prev[8][151] & 1'b1;
			partial_clause[8][152] 	= partial_clause_prev[8][152] & 1'b1;
			partial_clause[8][153] 	= partial_clause_prev[8][153] & 1'b1;
			partial_clause[8][154] 	= partial_clause_prev[8][154] & 1'b1;
			partial_clause[8][155] 	= partial_clause_prev[8][155] & 1'b1;
			partial_clause[8][156] 	= partial_clause_prev[8][156] & 1'b1;
			partial_clause[8][157] 	= partial_clause_prev[8][157] & 1'b1;
			partial_clause[8][158] 	= partial_clause_prev[8][158] & 1'b1;
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & 1'b1;
			partial_clause[8][161] 	= partial_clause_prev[8][161] & 1'b1;
			partial_clause[8][162] 	= partial_clause_prev[8][162] & 1'b1;
			partial_clause[8][163] 	= partial_clause_prev[8][163] & 1'b1;
			partial_clause[8][164] 	= partial_clause_prev[8][164] & 1'b1;
			partial_clause[8][165] 	= partial_clause_prev[8][165] & 1'b1;
			partial_clause[8][166] 	= partial_clause_prev[8][166] & 1'b1;
			partial_clause[8][167] 	= partial_clause_prev[8][167] & 1'b1;
			partial_clause[8][168] 	= partial_clause_prev[8][168] & 1'b1;
			partial_clause[8][169] 	= partial_clause_prev[8][169] & 1'b1;
			partial_clause[8][170] 	= partial_clause_prev[8][170] & x[34];
			partial_clause[8][171] 	= partial_clause_prev[8][171] & x[37];
			partial_clause[8][172] 	= partial_clause_prev[8][172] & 1'b1;
			partial_clause[8][173] 	= partial_clause_prev[8][173] & x[34];
			partial_clause[8][174] 	= partial_clause_prev[8][174] & 1'b1;
			partial_clause[8][175] 	= partial_clause_prev[8][175] & x[39];
			partial_clause[8][176] 	= partial_clause_prev[8][176] & 1'b1;
			partial_clause[8][177] 	= partial_clause_prev[8][177] & 1'b1;
			partial_clause[8][178] 	= partial_clause_prev[8][178] & 1'b1;
			partial_clause[8][179] 	= partial_clause_prev[8][179] & 1'b1;
			partial_clause[8][180] 	= partial_clause_prev[8][180] & 1'b1;
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & 1'b1;
			partial_clause[8][183] 	= partial_clause_prev[8][183] & 1'b1;
			partial_clause[8][184] 	= partial_clause_prev[8][184] & x[37];
			partial_clause[8][185] 	= partial_clause_prev[8][185] & 1'b1;
			partial_clause[8][186] 	= partial_clause_prev[8][186] & 1'b1;
			partial_clause[8][187] 	= partial_clause_prev[8][187] & 1'b1;
			partial_clause[8][188] 	= partial_clause_prev[8][188] & 1'b1;
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & 1'b1;
			partial_clause[8][191] 	= partial_clause_prev[8][191] & 1'b1;
			partial_clause[8][192] 	= partial_clause_prev[8][192] & 1'b1;
			partial_clause[8][193] 	= partial_clause_prev[8][193] & 1'b1;
			partial_clause[8][194] 	= partial_clause_prev[8][194] & 1'b1;
			partial_clause[8][195] 	= partial_clause_prev[8][195] & 1'b1;
			partial_clause[8][196] 	= partial_clause_prev[8][196] & 1'b1;
			partial_clause[8][197] 	= partial_clause_prev[8][197] & 1'b1;
			partial_clause[8][198] 	= partial_clause_prev[8][198] & 1'b1;
			partial_clause[8][199] 	= partial_clause_prev[8][199] & x[35];
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & x[4];
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & 1'b1;
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & x[39];
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & x[51];
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & x[41];
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
			partial_clause[9][100] 	= partial_clause_prev[9][100] & 1'b1;
			partial_clause[9][101] 	= partial_clause_prev[9][101] & 1'b1;
			partial_clause[9][102] 	= partial_clause_prev[9][102] & 1'b1;
			partial_clause[9][103] 	= partial_clause_prev[9][103] & 1'b1;
			partial_clause[9][104] 	= partial_clause_prev[9][104] & 1'b1;
			partial_clause[9][105] 	= partial_clause_prev[9][105] & 1'b1;
			partial_clause[9][106] 	= partial_clause_prev[9][106] & 1'b1;
			partial_clause[9][107] 	= partial_clause_prev[9][107] & 1'b1;
			partial_clause[9][108] 	= partial_clause_prev[9][108] & x[59];
			partial_clause[9][109] 	= partial_clause_prev[9][109] & 1'b1;
			partial_clause[9][110] 	= partial_clause_prev[9][110] & 1'b1;
			partial_clause[9][111] 	= partial_clause_prev[9][111] & 1'b1;
			partial_clause[9][112] 	= partial_clause_prev[9][112] & 1'b1;
			partial_clause[9][113] 	= partial_clause_prev[9][113] & 1'b1;
			partial_clause[9][114] 	= partial_clause_prev[9][114] & 1'b1;
			partial_clause[9][115] 	= partial_clause_prev[9][115] & 1'b1;
			partial_clause[9][116] 	= partial_clause_prev[9][116] & 1'b1;
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & 1'b1;
			partial_clause[9][119] 	= partial_clause_prev[9][119] & 1'b1;
			partial_clause[9][120] 	= partial_clause_prev[9][120] & 1'b1;
			partial_clause[9][121] 	= partial_clause_prev[9][121] & 1'b1;
			partial_clause[9][122] 	= partial_clause_prev[9][122] & 1'b1;
			partial_clause[9][123] 	= partial_clause_prev[9][123] & 1'b1;
			partial_clause[9][124] 	= partial_clause_prev[9][124] & 1'b1;
			partial_clause[9][125] 	= partial_clause_prev[9][125] & 1'b1;
			partial_clause[9][126] 	= partial_clause_prev[9][126] & 1'b1;
			partial_clause[9][127] 	= partial_clause_prev[9][127] & x[34];
			partial_clause[9][128] 	= partial_clause_prev[9][128] & x[63];
			partial_clause[9][129] 	= partial_clause_prev[9][129] & 1'b1;
			partial_clause[9][130] 	= partial_clause_prev[9][130] & 1'b1;
			partial_clause[9][131] 	= partial_clause_prev[9][131] & 1'b1;
			partial_clause[9][132] 	= partial_clause_prev[9][132] & 1'b1;
			partial_clause[9][133] 	= partial_clause_prev[9][133] & 1'b1;
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & 1'b1;
			partial_clause[9][138] 	= partial_clause_prev[9][138] & 1'b1;
			partial_clause[9][139] 	= partial_clause_prev[9][139] & 1'b1;
			partial_clause[9][140] 	= partial_clause_prev[9][140] & 1'b1;
			partial_clause[9][141] 	= partial_clause_prev[9][141] & 1'b1;
			partial_clause[9][142] 	= partial_clause_prev[9][142] & x[37];
			partial_clause[9][143] 	= partial_clause_prev[9][143] & 1'b1;
			partial_clause[9][144] 	= partial_clause_prev[9][144] & 1'b1;
			partial_clause[9][145] 	= partial_clause_prev[9][145] & 1'b1;
			partial_clause[9][146] 	= partial_clause_prev[9][146] & 1'b1;
			partial_clause[9][147] 	= partial_clause_prev[9][147] & 1'b1;
			partial_clause[9][148] 	= partial_clause_prev[9][148] & 1'b1;
			partial_clause[9][149] 	= partial_clause_prev[9][149] & ~x[25];
			partial_clause[9][150] 	= partial_clause_prev[9][150] & 1'b1;
			partial_clause[9][151] 	= partial_clause_prev[9][151] & 1'b1;
			partial_clause[9][152] 	= partial_clause_prev[9][152] & 1'b1;
			partial_clause[9][153] 	= partial_clause_prev[9][153] & 1'b1;
			partial_clause[9][154] 	= partial_clause_prev[9][154] & 1'b1;
			partial_clause[9][155] 	= partial_clause_prev[9][155] & 1'b1;
			partial_clause[9][156] 	= partial_clause_prev[9][156] & 1'b1;
			partial_clause[9][157] 	= partial_clause_prev[9][157] & 1'b1;
			partial_clause[9][158] 	= partial_clause_prev[9][158] & 1'b1;
			partial_clause[9][159] 	= partial_clause_prev[9][159] & x[62];
			partial_clause[9][160] 	= partial_clause_prev[9][160] & 1'b1;
			partial_clause[9][161] 	= partial_clause_prev[9][161] & 1'b1;
			partial_clause[9][162] 	= partial_clause_prev[9][162] & 1'b1;
			partial_clause[9][163] 	= partial_clause_prev[9][163] & 1'b1;
			partial_clause[9][164] 	= partial_clause_prev[9][164] & 1'b1;
			partial_clause[9][165] 	= partial_clause_prev[9][165] & 1'b1;
			partial_clause[9][166] 	= partial_clause_prev[9][166] & 1'b1;
			partial_clause[9][167] 	= partial_clause_prev[9][167] & 1'b1;
			partial_clause[9][168] 	= partial_clause_prev[9][168] & 1'b1;
			partial_clause[9][169] 	= partial_clause_prev[9][169] & 1'b1;
			partial_clause[9][170] 	= partial_clause_prev[9][170] & 1'b1;
			partial_clause[9][171] 	= partial_clause_prev[9][171] & 1'b1;
			partial_clause[9][172] 	= partial_clause_prev[9][172] & 1'b1;
			partial_clause[9][173] 	= partial_clause_prev[9][173] & 1'b1;
			partial_clause[9][174] 	= partial_clause_prev[9][174] & 1'b1;
			partial_clause[9][175] 	= partial_clause_prev[9][175] & 1'b1;
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & 1'b1;
			partial_clause[9][178] 	= partial_clause_prev[9][178] & 1'b1;
			partial_clause[9][179] 	= partial_clause_prev[9][179] & 1'b1;
			partial_clause[9][180] 	= partial_clause_prev[9][180] & 1'b1;
			partial_clause[9][181] 	= partial_clause_prev[9][181] & x[63];
			partial_clause[9][182] 	= partial_clause_prev[9][182] & ~x[51];
			partial_clause[9][183] 	= partial_clause_prev[9][183] & 1'b1;
			partial_clause[9][184] 	= partial_clause_prev[9][184] & 1'b1;
			partial_clause[9][185] 	= partial_clause_prev[9][185] & 1'b1;
			partial_clause[9][186] 	= partial_clause_prev[9][186] & x[61];
			partial_clause[9][187] 	= partial_clause_prev[9][187] & ~x[48];
			partial_clause[9][188] 	= partial_clause_prev[9][188] & 1'b1;
			partial_clause[9][189] 	= partial_clause_prev[9][189] & 1'b1;
			partial_clause[9][190] 	= partial_clause_prev[9][190] & 1'b1;
			partial_clause[9][191] 	= partial_clause_prev[9][191] & 1'b1;
			partial_clause[9][192] 	= partial_clause_prev[9][192] & 1'b1;
			partial_clause[9][193] 	= partial_clause_prev[9][193] & 1'b1;
			partial_clause[9][194] 	= partial_clause_prev[9][194] & 1'b1;
			partial_clause[9][195] 	= partial_clause_prev[9][195] & 1'b1;
			partial_clause[9][196] 	= partial_clause_prev[9][196] & 1'b1;
			partial_clause[9][197] 	= partial_clause_prev[9][197] & 1'b1;
			partial_clause[9][198] 	= partial_clause_prev[9][198] & 1'b1;
			partial_clause[9][199] 	= partial_clause_prev[9][199] & 1'b1;
		end
	end
endmodule


module HCB_2 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & ~x[23];
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & ~x[23];
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & x[13];
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & ~x[6];
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & ~x[13] & x[55];
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & ~x[50];
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & x[53];
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			partial_clause[0][100] 	= partial_clause_prev[0][100] & 1'b1;
			partial_clause[0][101] 	= partial_clause_prev[0][101] & 1'b1;
			partial_clause[0][102] 	= partial_clause_prev[0][102] & ~x[6];
			partial_clause[0][103] 	= partial_clause_prev[0][103] & 1'b1;
			partial_clause[0][104] 	= partial_clause_prev[0][104] & 1'b1;
			partial_clause[0][105] 	= partial_clause_prev[0][105] & 1'b1;
			partial_clause[0][106] 	= partial_clause_prev[0][106] & 1'b1;
			partial_clause[0][107] 	= partial_clause_prev[0][107] & 1'b1;
			partial_clause[0][108] 	= partial_clause_prev[0][108] & ~x[25] & ~x[27];
			partial_clause[0][109] 	= partial_clause_prev[0][109] & 1'b1;
			partial_clause[0][110] 	= partial_clause_prev[0][110] & 1'b1;
			partial_clause[0][111] 	= partial_clause_prev[0][111] & 1'b1;
			partial_clause[0][112] 	= partial_clause_prev[0][112] & 1'b1;
			partial_clause[0][113] 	= partial_clause_prev[0][113] & 1'b1;
			partial_clause[0][114] 	= partial_clause_prev[0][114] & 1'b1;
			partial_clause[0][115] 	= partial_clause_prev[0][115] & 1'b1;
			partial_clause[0][116] 	= partial_clause_prev[0][116] & 1'b1;
			partial_clause[0][117] 	= partial_clause_prev[0][117] & 1'b1;
			partial_clause[0][118] 	= partial_clause_prev[0][118] & 1'b1;
			partial_clause[0][119] 	= partial_clause_prev[0][119] & 1'b1;
			partial_clause[0][120] 	= partial_clause_prev[0][120] & 1'b1;
			partial_clause[0][121] 	= partial_clause_prev[0][121] & 1'b1;
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & 1'b1;
			partial_clause[0][124] 	= partial_clause_prev[0][124] & 1'b1;
			partial_clause[0][125] 	= partial_clause_prev[0][125] & 1'b1;
			partial_clause[0][126] 	= partial_clause_prev[0][126] & 1'b1;
			partial_clause[0][127] 	= partial_clause_prev[0][127] & 1'b1;
			partial_clause[0][128] 	= partial_clause_prev[0][128] & ~x[26] & ~x[57];
			partial_clause[0][129] 	= partial_clause_prev[0][129] & 1'b1;
			partial_clause[0][130] 	= partial_clause_prev[0][130] & 1'b1;
			partial_clause[0][131] 	= partial_clause_prev[0][131] & 1'b1;
			partial_clause[0][132] 	= partial_clause_prev[0][132] & 1'b1;
			partial_clause[0][133] 	= partial_clause_prev[0][133] & 1'b1;
			partial_clause[0][134] 	= partial_clause_prev[0][134] & 1'b1;
			partial_clause[0][135] 	= partial_clause_prev[0][135] & 1'b1;
			partial_clause[0][136] 	= partial_clause_prev[0][136] & 1'b1;
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & ~x[0] & ~x[25];
			partial_clause[0][139] 	= partial_clause_prev[0][139] & 1'b1;
			partial_clause[0][140] 	= partial_clause_prev[0][140] & x[21];
			partial_clause[0][141] 	= partial_clause_prev[0][141] & 1'b1;
			partial_clause[0][142] 	= partial_clause_prev[0][142] & 1'b1;
			partial_clause[0][143] 	= partial_clause_prev[0][143] & 1'b1;
			partial_clause[0][144] 	= partial_clause_prev[0][144] & 1'b1;
			partial_clause[0][145] 	= partial_clause_prev[0][145] & 1'b1;
			partial_clause[0][146] 	= partial_clause_prev[0][146] & 1'b1;
			partial_clause[0][147] 	= partial_clause_prev[0][147] & 1'b1;
			partial_clause[0][148] 	= partial_clause_prev[0][148] & 1'b1;
			partial_clause[0][149] 	= partial_clause_prev[0][149] & 1'b1;
			partial_clause[0][150] 	= partial_clause_prev[0][150] & 1'b1;
			partial_clause[0][151] 	= partial_clause_prev[0][151] & 1'b1;
			partial_clause[0][152] 	= partial_clause_prev[0][152] & 1'b1;
			partial_clause[0][153] 	= partial_clause_prev[0][153] & 1'b1;
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & 1'b1;
			partial_clause[0][156] 	= partial_clause_prev[0][156] & 1'b1;
			partial_clause[0][157] 	= partial_clause_prev[0][157] & 1'b1;
			partial_clause[0][158] 	= partial_clause_prev[0][158] & 1'b1;
			partial_clause[0][159] 	= partial_clause_prev[0][159] & 1'b1;
			partial_clause[0][160] 	= partial_clause_prev[0][160] & 1'b1;
			partial_clause[0][161] 	= partial_clause_prev[0][161] & 1'b1;
			partial_clause[0][162] 	= partial_clause_prev[0][162] & 1'b1;
			partial_clause[0][163] 	= partial_clause_prev[0][163] & 1'b1;
			partial_clause[0][164] 	= partial_clause_prev[0][164] & 1'b1;
			partial_clause[0][165] 	= partial_clause_prev[0][165] & 1'b1;
			partial_clause[0][166] 	= partial_clause_prev[0][166] & 1'b1;
			partial_clause[0][167] 	= partial_clause_prev[0][167] & 1'b1;
			partial_clause[0][168] 	= partial_clause_prev[0][168] & 1'b1;
			partial_clause[0][169] 	= partial_clause_prev[0][169] & 1'b1;
			partial_clause[0][170] 	= partial_clause_prev[0][170] & 1'b1;
			partial_clause[0][171] 	= partial_clause_prev[0][171] & 1'b1;
			partial_clause[0][172] 	= partial_clause_prev[0][172] & 1'b1;
			partial_clause[0][173] 	= partial_clause_prev[0][173] & 1'b1;
			partial_clause[0][174] 	= partial_clause_prev[0][174] & 1'b1;
			partial_clause[0][175] 	= partial_clause_prev[0][175] & 1'b1;
			partial_clause[0][176] 	= partial_clause_prev[0][176] & 1'b1;
			partial_clause[0][177] 	= partial_clause_prev[0][177] & 1'b1;
			partial_clause[0][178] 	= partial_clause_prev[0][178] & 1'b1;
			partial_clause[0][179] 	= partial_clause_prev[0][179] & 1'b1;
			partial_clause[0][180] 	= partial_clause_prev[0][180] & 1'b1;
			partial_clause[0][181] 	= partial_clause_prev[0][181] & 1'b1;
			partial_clause[0][182] 	= partial_clause_prev[0][182] & 1'b1;
			partial_clause[0][183] 	= partial_clause_prev[0][183] & 1'b1;
			partial_clause[0][184] 	= partial_clause_prev[0][184] & 1'b1;
			partial_clause[0][185] 	= partial_clause_prev[0][185] & x[48];
			partial_clause[0][186] 	= partial_clause_prev[0][186] & 1'b1;
			partial_clause[0][187] 	= partial_clause_prev[0][187] & 1'b1;
			partial_clause[0][188] 	= partial_clause_prev[0][188] & 1'b1;
			partial_clause[0][189] 	= partial_clause_prev[0][189] & 1'b1;
			partial_clause[0][190] 	= partial_clause_prev[0][190] & 1'b1;
			partial_clause[0][191] 	= partial_clause_prev[0][191] & 1'b1;
			partial_clause[0][192] 	= partial_clause_prev[0][192] & 1'b1;
			partial_clause[0][193] 	= partial_clause_prev[0][193] & 1'b1;
			partial_clause[0][194] 	= partial_clause_prev[0][194] & 1'b1;
			partial_clause[0][195] 	= partial_clause_prev[0][195] & 1'b1;
			partial_clause[0][196] 	= partial_clause_prev[0][196] & ~x[25] & ~x[30] & ~x[55];
			partial_clause[0][197] 	= partial_clause_prev[0][197] & 1'b1;
			partial_clause[0][198] 	= partial_clause_prev[0][198] & 1'b1;
			partial_clause[0][199] 	= partial_clause_prev[0][199] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[53];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & x[26] & ~x[49];
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & x[15];
			partial_clause[1][15] 	= partial_clause_prev[1][15] & ~x[49];
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & x[38];
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & ~x[49] & ~x[51];
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & x[15];
			partial_clause[1][38] 	= partial_clause_prev[1][38] & x[45];
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & x[16];
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & ~x[58];
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & x[33];
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & ~x[26];
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & ~x[54];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & ~x[27] & ~x[28];
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & ~x[49];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & ~x[60];
			partial_clause[1][78] 	= partial_clause_prev[1][78] & ~x[54];
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & ~x[25];
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			partial_clause[1][100] 	= partial_clause_prev[1][100] & 1'b1;
			partial_clause[1][101] 	= partial_clause_prev[1][101] & x[54] & x[57];
			partial_clause[1][102] 	= partial_clause_prev[1][102] & 1'b1;
			partial_clause[1][103] 	= partial_clause_prev[1][103] & 1'b1;
			partial_clause[1][104] 	= partial_clause_prev[1][104] & 1'b1;
			partial_clause[1][105] 	= partial_clause_prev[1][105] & 1'b1;
			partial_clause[1][106] 	= partial_clause_prev[1][106] & 1'b1;
			partial_clause[1][107] 	= partial_clause_prev[1][107] & 1'b1;
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & x[54] & x[55];
			partial_clause[1][110] 	= partial_clause_prev[1][110] & ~x[23];
			partial_clause[1][111] 	= partial_clause_prev[1][111] & 1'b1;
			partial_clause[1][112] 	= partial_clause_prev[1][112] & 1'b1;
			partial_clause[1][113] 	= partial_clause_prev[1][113] & 1'b1;
			partial_clause[1][114] 	= partial_clause_prev[1][114] & 1'b1;
			partial_clause[1][115] 	= partial_clause_prev[1][115] & 1'b1;
			partial_clause[1][116] 	= partial_clause_prev[1][116] & 1'b1;
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & 1'b1;
			partial_clause[1][119] 	= partial_clause_prev[1][119] & 1'b1;
			partial_clause[1][120] 	= partial_clause_prev[1][120] & 1'b1;
			partial_clause[1][121] 	= partial_clause_prev[1][121] & 1'b1;
			partial_clause[1][122] 	= partial_clause_prev[1][122] & 1'b1;
			partial_clause[1][123] 	= partial_clause_prev[1][123] & 1'b1;
			partial_clause[1][124] 	= partial_clause_prev[1][124] & x[51];
			partial_clause[1][125] 	= partial_clause_prev[1][125] & 1'b1;
			partial_clause[1][126] 	= partial_clause_prev[1][126] & 1'b1;
			partial_clause[1][127] 	= partial_clause_prev[1][127] & 1'b1;
			partial_clause[1][128] 	= partial_clause_prev[1][128] & ~x[16];
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & ~x[30] & ~x[31] & ~x[40];
			partial_clause[1][131] 	= partial_clause_prev[1][131] & 1'b1;
			partial_clause[1][132] 	= partial_clause_prev[1][132] & 1'b1;
			partial_clause[1][133] 	= partial_clause_prev[1][133] & 1'b1;
			partial_clause[1][134] 	= partial_clause_prev[1][134] & 1'b1;
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & 1'b1;
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & 1'b1;
			partial_clause[1][139] 	= partial_clause_prev[1][139] & 1'b1;
			partial_clause[1][140] 	= partial_clause_prev[1][140] & 1'b1;
			partial_clause[1][141] 	= partial_clause_prev[1][141] & 1'b1;
			partial_clause[1][142] 	= partial_clause_prev[1][142] & 1'b1;
			partial_clause[1][143] 	= partial_clause_prev[1][143] & 1'b1;
			partial_clause[1][144] 	= partial_clause_prev[1][144] & 1'b1;
			partial_clause[1][145] 	= partial_clause_prev[1][145] & 1'b1;
			partial_clause[1][146] 	= partial_clause_prev[1][146] & x[24];
			partial_clause[1][147] 	= partial_clause_prev[1][147] & x[52];
			partial_clause[1][148] 	= partial_clause_prev[1][148] & 1'b1;
			partial_clause[1][149] 	= partial_clause_prev[1][149] & 1'b1;
			partial_clause[1][150] 	= partial_clause_prev[1][150] & 1'b1;
			partial_clause[1][151] 	= partial_clause_prev[1][151] & x[49];
			partial_clause[1][152] 	= partial_clause_prev[1][152] & 1'b1;
			partial_clause[1][153] 	= partial_clause_prev[1][153] & 1'b1;
			partial_clause[1][154] 	= partial_clause_prev[1][154] & 1'b1;
			partial_clause[1][155] 	= partial_clause_prev[1][155] & 1'b1;
			partial_clause[1][156] 	= partial_clause_prev[1][156] & 1'b1;
			partial_clause[1][157] 	= partial_clause_prev[1][157] & 1'b1;
			partial_clause[1][158] 	= partial_clause_prev[1][158] & 1'b1;
			partial_clause[1][159] 	= partial_clause_prev[1][159] & ~x[0] & ~x[27];
			partial_clause[1][160] 	= partial_clause_prev[1][160] & 1'b1;
			partial_clause[1][161] 	= partial_clause_prev[1][161] & 1'b1;
			partial_clause[1][162] 	= partial_clause_prev[1][162] & 1'b1;
			partial_clause[1][163] 	= partial_clause_prev[1][163] & ~x[29];
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & 1'b1;
			partial_clause[1][166] 	= partial_clause_prev[1][166] & 1'b1;
			partial_clause[1][167] 	= partial_clause_prev[1][167] & 1'b1;
			partial_clause[1][168] 	= partial_clause_prev[1][168] & 1'b1;
			partial_clause[1][169] 	= partial_clause_prev[1][169] & 1'b1;
			partial_clause[1][170] 	= partial_clause_prev[1][170] & x[20];
			partial_clause[1][171] 	= partial_clause_prev[1][171] & 1'b1;
			partial_clause[1][172] 	= partial_clause_prev[1][172] & 1'b1;
			partial_clause[1][173] 	= partial_clause_prev[1][173] & 1'b1;
			partial_clause[1][174] 	= partial_clause_prev[1][174] & 1'b1;
			partial_clause[1][175] 	= partial_clause_prev[1][175] & 1'b1;
			partial_clause[1][176] 	= partial_clause_prev[1][176] & 1'b1;
			partial_clause[1][177] 	= partial_clause_prev[1][177] & ~x[27];
			partial_clause[1][178] 	= partial_clause_prev[1][178] & 1'b1;
			partial_clause[1][179] 	= partial_clause_prev[1][179] & 1'b1;
			partial_clause[1][180] 	= partial_clause_prev[1][180] & 1'b1;
			partial_clause[1][181] 	= partial_clause_prev[1][181] & 1'b1;
			partial_clause[1][182] 	= partial_clause_prev[1][182] & 1'b1;
			partial_clause[1][183] 	= partial_clause_prev[1][183] & 1'b1;
			partial_clause[1][184] 	= partial_clause_prev[1][184] & ~x[31];
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & 1'b1;
			partial_clause[1][187] 	= partial_clause_prev[1][187] & 1'b1;
			partial_clause[1][188] 	= partial_clause_prev[1][188] & x[23];
			partial_clause[1][189] 	= partial_clause_prev[1][189] & 1'b1;
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & 1'b1;
			partial_clause[1][192] 	= partial_clause_prev[1][192] & 1'b1;
			partial_clause[1][193] 	= partial_clause_prev[1][193] & 1'b1;
			partial_clause[1][194] 	= partial_clause_prev[1][194] & 1'b1;
			partial_clause[1][195] 	= partial_clause_prev[1][195] & 1'b1;
			partial_clause[1][196] 	= partial_clause_prev[1][196] & x[25];
			partial_clause[1][197] 	= partial_clause_prev[1][197] & 1'b1;
			partial_clause[1][198] 	= partial_clause_prev[1][198] & 1'b1;
			partial_clause[1][199] 	= partial_clause_prev[1][199] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & x[24];
			partial_clause[2][2] 	= partial_clause_prev[2][2] & x[54];
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & x[27];
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & x[27];
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & x[1];
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & x[28];
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & x[0];
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & x[27];
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & x[25];
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & x[54];
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & ~x[9];
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & x[23];
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & 1'b1;
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & x[55];
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			partial_clause[2][100] 	= partial_clause_prev[2][100] & 1'b1;
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & 1'b1;
			partial_clause[2][103] 	= partial_clause_prev[2][103] & 1'b1;
			partial_clause[2][104] 	= partial_clause_prev[2][104] & 1'b1;
			partial_clause[2][105] 	= partial_clause_prev[2][105] & 1'b1;
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & 1'b1;
			partial_clause[2][108] 	= partial_clause_prev[2][108] & 1'b1;
			partial_clause[2][109] 	= partial_clause_prev[2][109] & 1'b1;
			partial_clause[2][110] 	= partial_clause_prev[2][110] & 1'b1;
			partial_clause[2][111] 	= partial_clause_prev[2][111] & 1'b1;
			partial_clause[2][112] 	= partial_clause_prev[2][112] & 1'b1;
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & 1'b1;
			partial_clause[2][115] 	= partial_clause_prev[2][115] & 1'b1;
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & 1'b1;
			partial_clause[2][118] 	= partial_clause_prev[2][118] & 1'b1;
			partial_clause[2][119] 	= partial_clause_prev[2][119] & 1'b1;
			partial_clause[2][120] 	= partial_clause_prev[2][120] & 1'b1;
			partial_clause[2][121] 	= partial_clause_prev[2][121] & 1'b1;
			partial_clause[2][122] 	= partial_clause_prev[2][122] & 1'b1;
			partial_clause[2][123] 	= partial_clause_prev[2][123] & 1'b1;
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & 1'b1;
			partial_clause[2][126] 	= partial_clause_prev[2][126] & 1'b1;
			partial_clause[2][127] 	= partial_clause_prev[2][127] & 1'b1;
			partial_clause[2][128] 	= partial_clause_prev[2][128] & 1'b1;
			partial_clause[2][129] 	= partial_clause_prev[2][129] & 1'b1;
			partial_clause[2][130] 	= partial_clause_prev[2][130] & 1'b1;
			partial_clause[2][131] 	= partial_clause_prev[2][131] & 1'b1;
			partial_clause[2][132] 	= partial_clause_prev[2][132] & 1'b1;
			partial_clause[2][133] 	= partial_clause_prev[2][133] & 1'b1;
			partial_clause[2][134] 	= partial_clause_prev[2][134] & 1'b1;
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & 1'b1;
			partial_clause[2][137] 	= partial_clause_prev[2][137] & 1'b1;
			partial_clause[2][138] 	= partial_clause_prev[2][138] & 1'b1;
			partial_clause[2][139] 	= partial_clause_prev[2][139] & 1'b1;
			partial_clause[2][140] 	= partial_clause_prev[2][140] & 1'b1;
			partial_clause[2][141] 	= partial_clause_prev[2][141] & 1'b1;
			partial_clause[2][142] 	= partial_clause_prev[2][142] & 1'b1;
			partial_clause[2][143] 	= partial_clause_prev[2][143] & 1'b1;
			partial_clause[2][144] 	= partial_clause_prev[2][144] & 1'b1;
			partial_clause[2][145] 	= partial_clause_prev[2][145] & 1'b1;
			partial_clause[2][146] 	= partial_clause_prev[2][146] & 1'b1;
			partial_clause[2][147] 	= partial_clause_prev[2][147] & 1'b1;
			partial_clause[2][148] 	= partial_clause_prev[2][148] & 1'b1;
			partial_clause[2][149] 	= partial_clause_prev[2][149] & 1'b1;
			partial_clause[2][150] 	= partial_clause_prev[2][150] & 1'b1;
			partial_clause[2][151] 	= partial_clause_prev[2][151] & x[6];
			partial_clause[2][152] 	= partial_clause_prev[2][152] & 1'b1;
			partial_clause[2][153] 	= partial_clause_prev[2][153] & 1'b1;
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & 1'b1;
			partial_clause[2][156] 	= partial_clause_prev[2][156] & 1'b1;
			partial_clause[2][157] 	= partial_clause_prev[2][157] & 1'b1;
			partial_clause[2][158] 	= partial_clause_prev[2][158] & 1'b1;
			partial_clause[2][159] 	= partial_clause_prev[2][159] & 1'b1;
			partial_clause[2][160] 	= partial_clause_prev[2][160] & 1'b1;
			partial_clause[2][161] 	= partial_clause_prev[2][161] & 1'b1;
			partial_clause[2][162] 	= partial_clause_prev[2][162] & 1'b1;
			partial_clause[2][163] 	= partial_clause_prev[2][163] & 1'b1;
			partial_clause[2][164] 	= partial_clause_prev[2][164] & 1'b1;
			partial_clause[2][165] 	= partial_clause_prev[2][165] & 1'b1;
			partial_clause[2][166] 	= partial_clause_prev[2][166] & 1'b1;
			partial_clause[2][167] 	= partial_clause_prev[2][167] & 1'b1;
			partial_clause[2][168] 	= partial_clause_prev[2][168] & 1'b1;
			partial_clause[2][169] 	= partial_clause_prev[2][169] & 1'b1;
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & 1'b1;
			partial_clause[2][173] 	= partial_clause_prev[2][173] & 1'b1;
			partial_clause[2][174] 	= partial_clause_prev[2][174] & 1'b1;
			partial_clause[2][175] 	= partial_clause_prev[2][175] & 1'b1;
			partial_clause[2][176] 	= partial_clause_prev[2][176] & 1'b1;
			partial_clause[2][177] 	= partial_clause_prev[2][177] & ~x[26];
			partial_clause[2][178] 	= partial_clause_prev[2][178] & 1'b1;
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & 1'b1;
			partial_clause[2][181] 	= partial_clause_prev[2][181] & ~x[48];
			partial_clause[2][182] 	= partial_clause_prev[2][182] & 1'b1;
			partial_clause[2][183] 	= partial_clause_prev[2][183] & 1'b1;
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & 1'b1;
			partial_clause[2][186] 	= partial_clause_prev[2][186] & 1'b1;
			partial_clause[2][187] 	= partial_clause_prev[2][187] & 1'b1;
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & ~x[48];
			partial_clause[2][190] 	= partial_clause_prev[2][190] & 1'b1;
			partial_clause[2][191] 	= partial_clause_prev[2][191] & 1'b1;
			partial_clause[2][192] 	= partial_clause_prev[2][192] & 1'b1;
			partial_clause[2][193] 	= partial_clause_prev[2][193] & 1'b1;
			partial_clause[2][194] 	= partial_clause_prev[2][194] & 1'b1;
			partial_clause[2][195] 	= partial_clause_prev[2][195] & 1'b1;
			partial_clause[2][196] 	= partial_clause_prev[2][196] & 1'b1;
			partial_clause[2][197] 	= partial_clause_prev[2][197] & 1'b1;
			partial_clause[2][198] 	= partial_clause_prev[2][198] & 1'b1;
			partial_clause[2][199] 	= partial_clause_prev[2][199] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & x[49];
			partial_clause[3][2] 	= partial_clause_prev[3][2] & x[52];
			partial_clause[3][3] 	= partial_clause_prev[3][3] & x[53];
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & x[17];
			partial_clause[3][8] 	= partial_clause_prev[3][8] & x[18];
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & x[26];
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & x[24];
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & ~x[60];
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & x[26];
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & x[53];
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & x[51];
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & x[55];
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & x[11];
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & x[23];
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & ~x[27];
			partial_clause[3][63] 	= partial_clause_prev[3][63] & x[56];
			partial_clause[3][64] 	= partial_clause_prev[3][64] & x[45];
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[31];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & x[25];
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & x[10];
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & x[22];
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & x[27];
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & x[44];
			partial_clause[3][100] 	= partial_clause_prev[3][100] & 1'b1;
			partial_clause[3][101] 	= partial_clause_prev[3][101] & 1'b1;
			partial_clause[3][102] 	= partial_clause_prev[3][102] & 1'b1;
			partial_clause[3][103] 	= partial_clause_prev[3][103] & 1'b1;
			partial_clause[3][104] 	= partial_clause_prev[3][104] & 1'b1;
			partial_clause[3][105] 	= partial_clause_prev[3][105] & 1'b1;
			partial_clause[3][106] 	= partial_clause_prev[3][106] & 1'b1;
			partial_clause[3][107] 	= partial_clause_prev[3][107] & 1'b1;
			partial_clause[3][108] 	= partial_clause_prev[3][108] & 1'b1;
			partial_clause[3][109] 	= partial_clause_prev[3][109] & 1'b1;
			partial_clause[3][110] 	= partial_clause_prev[3][110] & 1'b1;
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & 1'b1;
			partial_clause[3][113] 	= partial_clause_prev[3][113] & ~x[50];
			partial_clause[3][114] 	= partial_clause_prev[3][114] & 1'b1;
			partial_clause[3][115] 	= partial_clause_prev[3][115] & 1'b1;
			partial_clause[3][116] 	= partial_clause_prev[3][116] & 1'b1;
			partial_clause[3][117] 	= partial_clause_prev[3][117] & 1'b1;
			partial_clause[3][118] 	= partial_clause_prev[3][118] & 1'b1;
			partial_clause[3][119] 	= partial_clause_prev[3][119] & 1'b1;
			partial_clause[3][120] 	= partial_clause_prev[3][120] & 1'b1;
			partial_clause[3][121] 	= partial_clause_prev[3][121] & 1'b1;
			partial_clause[3][122] 	= partial_clause_prev[3][122] & 1'b1;
			partial_clause[3][123] 	= partial_clause_prev[3][123] & 1'b1;
			partial_clause[3][124] 	= partial_clause_prev[3][124] & 1'b1;
			partial_clause[3][125] 	= partial_clause_prev[3][125] & 1'b1;
			partial_clause[3][126] 	= partial_clause_prev[3][126] & 1'b1;
			partial_clause[3][127] 	= partial_clause_prev[3][127] & 1'b1;
			partial_clause[3][128] 	= partial_clause_prev[3][128] & ~x[22];
			partial_clause[3][129] 	= partial_clause_prev[3][129] & 1'b1;
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & 1'b1;
			partial_clause[3][132] 	= partial_clause_prev[3][132] & 1'b1;
			partial_clause[3][133] 	= partial_clause_prev[3][133] & ~x[23] & ~x[56];
			partial_clause[3][134] 	= partial_clause_prev[3][134] & 1'b1;
			partial_clause[3][135] 	= partial_clause_prev[3][135] & 1'b1;
			partial_clause[3][136] 	= partial_clause_prev[3][136] & 1'b1;
			partial_clause[3][137] 	= partial_clause_prev[3][137] & 1'b1;
			partial_clause[3][138] 	= partial_clause_prev[3][138] & 1'b1;
			partial_clause[3][139] 	= partial_clause_prev[3][139] & 1'b1;
			partial_clause[3][140] 	= partial_clause_prev[3][140] & 1'b1;
			partial_clause[3][141] 	= partial_clause_prev[3][141] & 1'b1;
			partial_clause[3][142] 	= partial_clause_prev[3][142] & 1'b1;
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & 1'b1;
			partial_clause[3][145] 	= partial_clause_prev[3][145] & ~x[22] & ~x[50];
			partial_clause[3][146] 	= partial_clause_prev[3][146] & 1'b1;
			partial_clause[3][147] 	= partial_clause_prev[3][147] & 1'b1;
			partial_clause[3][148] 	= partial_clause_prev[3][148] & 1'b1;
			partial_clause[3][149] 	= partial_clause_prev[3][149] & 1'b1;
			partial_clause[3][150] 	= partial_clause_prev[3][150] & x[34];
			partial_clause[3][151] 	= partial_clause_prev[3][151] & 1'b1;
			partial_clause[3][152] 	= partial_clause_prev[3][152] & 1'b1;
			partial_clause[3][153] 	= partial_clause_prev[3][153] & 1'b1;
			partial_clause[3][154] 	= partial_clause_prev[3][154] & 1'b1;
			partial_clause[3][155] 	= partial_clause_prev[3][155] & 1'b1;
			partial_clause[3][156] 	= partial_clause_prev[3][156] & 1'b1;
			partial_clause[3][157] 	= partial_clause_prev[3][157] & 1'b1;
			partial_clause[3][158] 	= partial_clause_prev[3][158] & 1'b1;
			partial_clause[3][159] 	= partial_clause_prev[3][159] & 1'b1;
			partial_clause[3][160] 	= partial_clause_prev[3][160] & 1'b1;
			partial_clause[3][161] 	= partial_clause_prev[3][161] & 1'b1;
			partial_clause[3][162] 	= partial_clause_prev[3][162] & 1'b1;
			partial_clause[3][163] 	= partial_clause_prev[3][163] & 1'b1;
			partial_clause[3][164] 	= partial_clause_prev[3][164] & 1'b1;
			partial_clause[3][165] 	= partial_clause_prev[3][165] & x[35];
			partial_clause[3][166] 	= partial_clause_prev[3][166] & 1'b1;
			partial_clause[3][167] 	= partial_clause_prev[3][167] & 1'b1;
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & 1'b1;
			partial_clause[3][170] 	= partial_clause_prev[3][170] & 1'b1;
			partial_clause[3][171] 	= partial_clause_prev[3][171] & 1'b1;
			partial_clause[3][172] 	= partial_clause_prev[3][172] & 1'b1;
			partial_clause[3][173] 	= partial_clause_prev[3][173] & ~x[24] & ~x[51];
			partial_clause[3][174] 	= partial_clause_prev[3][174] & 1'b1;
			partial_clause[3][175] 	= partial_clause_prev[3][175] & 1'b1;
			partial_clause[3][176] 	= partial_clause_prev[3][176] & 1'b1;
			partial_clause[3][177] 	= partial_clause_prev[3][177] & ~x[49];
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & x[63];
			partial_clause[3][180] 	= partial_clause_prev[3][180] & ~x[49];
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & 1'b1;
			partial_clause[3][183] 	= partial_clause_prev[3][183] & 1'b1;
			partial_clause[3][184] 	= partial_clause_prev[3][184] & 1'b1;
			partial_clause[3][185] 	= partial_clause_prev[3][185] & 1'b1;
			partial_clause[3][186] 	= partial_clause_prev[3][186] & 1'b1;
			partial_clause[3][187] 	= partial_clause_prev[3][187] & 1'b1;
			partial_clause[3][188] 	= partial_clause_prev[3][188] & x[36];
			partial_clause[3][189] 	= partial_clause_prev[3][189] & 1'b1;
			partial_clause[3][190] 	= partial_clause_prev[3][190] & 1'b1;
			partial_clause[3][191] 	= partial_clause_prev[3][191] & 1'b1;
			partial_clause[3][192] 	= partial_clause_prev[3][192] & 1'b1;
			partial_clause[3][193] 	= partial_clause_prev[3][193] & 1'b1;
			partial_clause[3][194] 	= partial_clause_prev[3][194] & 1'b1;
			partial_clause[3][195] 	= partial_clause_prev[3][195] & 1'b1;
			partial_clause[3][196] 	= partial_clause_prev[3][196] & 1'b1;
			partial_clause[3][197] 	= partial_clause_prev[3][197] & 1'b1;
			partial_clause[3][198] 	= partial_clause_prev[3][198] & 1'b1;
			partial_clause[3][199] 	= partial_clause_prev[3][199] & ~x[22] & ~x[24];
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & ~x[55];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & ~x[53];
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & ~x[26];
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & ~x[0] & ~x[58];
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & x[63];
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & x[62];
			partial_clause[4][26] 	= partial_clause_prev[4][26] & x[63];
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[55];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & ~x[50];
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & ~x[27];
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & x[10];
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[54];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & ~x[54];
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & ~x[53];
			partial_clause[4][53] 	= partial_clause_prev[4][53] & ~x[28];
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & ~x[54];
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & x[11];
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & ~x[54];
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & ~x[28] & ~x[55];
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & x[41];
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			partial_clause[4][100] 	= partial_clause_prev[4][100] & 1'b1;
			partial_clause[4][101] 	= partial_clause_prev[4][101] & 1'b1;
			partial_clause[4][102] 	= partial_clause_prev[4][102] & 1'b1;
			partial_clause[4][103] 	= partial_clause_prev[4][103] & 1'b1;
			partial_clause[4][104] 	= partial_clause_prev[4][104] & 1'b1;
			partial_clause[4][105] 	= partial_clause_prev[4][105] & x[51];
			partial_clause[4][106] 	= partial_clause_prev[4][106] & 1'b1;
			partial_clause[4][107] 	= partial_clause_prev[4][107] & 1'b1;
			partial_clause[4][108] 	= partial_clause_prev[4][108] & 1'b1;
			partial_clause[4][109] 	= partial_clause_prev[4][109] & ~x[26];
			partial_clause[4][110] 	= partial_clause_prev[4][110] & 1'b1;
			partial_clause[4][111] 	= partial_clause_prev[4][111] & 1'b1;
			partial_clause[4][112] 	= partial_clause_prev[4][112] & 1'b1;
			partial_clause[4][113] 	= partial_clause_prev[4][113] & 1'b1;
			partial_clause[4][114] 	= partial_clause_prev[4][114] & 1'b1;
			partial_clause[4][115] 	= partial_clause_prev[4][115] & 1'b1;
			partial_clause[4][116] 	= partial_clause_prev[4][116] & 1'b1;
			partial_clause[4][117] 	= partial_clause_prev[4][117] & 1'b1;
			partial_clause[4][118] 	= partial_clause_prev[4][118] & 1'b1;
			partial_clause[4][119] 	= partial_clause_prev[4][119] & 1'b1;
			partial_clause[4][120] 	= partial_clause_prev[4][120] & 1'b1;
			partial_clause[4][121] 	= partial_clause_prev[4][121] & 1'b1;
			partial_clause[4][122] 	= partial_clause_prev[4][122] & 1'b1;
			partial_clause[4][123] 	= partial_clause_prev[4][123] & 1'b1;
			partial_clause[4][124] 	= partial_clause_prev[4][124] & 1'b1;
			partial_clause[4][125] 	= partial_clause_prev[4][125] & 1'b1;
			partial_clause[4][126] 	= partial_clause_prev[4][126] & 1'b1;
			partial_clause[4][127] 	= partial_clause_prev[4][127] & 1'b1;
			partial_clause[4][128] 	= partial_clause_prev[4][128] & 1'b1;
			partial_clause[4][129] 	= partial_clause_prev[4][129] & 1'b1;
			partial_clause[4][130] 	= partial_clause_prev[4][130] & 1'b1;
			partial_clause[4][131] 	= partial_clause_prev[4][131] & 1'b1;
			partial_clause[4][132] 	= partial_clause_prev[4][132] & 1'b1;
			partial_clause[4][133] 	= partial_clause_prev[4][133] & 1'b1;
			partial_clause[4][134] 	= partial_clause_prev[4][134] & 1'b1;
			partial_clause[4][135] 	= partial_clause_prev[4][135] & 1'b1;
			partial_clause[4][136] 	= partial_clause_prev[4][136] & 1'b1;
			partial_clause[4][137] 	= partial_clause_prev[4][137] & 1'b1;
			partial_clause[4][138] 	= partial_clause_prev[4][138] & 1'b1;
			partial_clause[4][139] 	= partial_clause_prev[4][139] & 1'b1;
			partial_clause[4][140] 	= partial_clause_prev[4][140] & 1'b1;
			partial_clause[4][141] 	= partial_clause_prev[4][141] & 1'b1;
			partial_clause[4][142] 	= partial_clause_prev[4][142] & 1'b1;
			partial_clause[4][143] 	= partial_clause_prev[4][143] & ~x[30];
			partial_clause[4][144] 	= partial_clause_prev[4][144] & 1'b1;
			partial_clause[4][145] 	= partial_clause_prev[4][145] & 1'b1;
			partial_clause[4][146] 	= partial_clause_prev[4][146] & x[30];
			partial_clause[4][147] 	= partial_clause_prev[4][147] & 1'b1;
			partial_clause[4][148] 	= partial_clause_prev[4][148] & x[52];
			partial_clause[4][149] 	= partial_clause_prev[4][149] & 1'b1;
			partial_clause[4][150] 	= partial_clause_prev[4][150] & 1'b1;
			partial_clause[4][151] 	= partial_clause_prev[4][151] & x[55];
			partial_clause[4][152] 	= partial_clause_prev[4][152] & 1'b1;
			partial_clause[4][153] 	= partial_clause_prev[4][153] & 1'b1;
			partial_clause[4][154] 	= partial_clause_prev[4][154] & x[25];
			partial_clause[4][155] 	= partial_clause_prev[4][155] & 1'b1;
			partial_clause[4][156] 	= partial_clause_prev[4][156] & 1'b1;
			partial_clause[4][157] 	= partial_clause_prev[4][157] & ~x[26] & ~x[28];
			partial_clause[4][158] 	= partial_clause_prev[4][158] & 1'b1;
			partial_clause[4][159] 	= partial_clause_prev[4][159] & 1'b1;
			partial_clause[4][160] 	= partial_clause_prev[4][160] & ~x[27];
			partial_clause[4][161] 	= partial_clause_prev[4][161] & 1'b1;
			partial_clause[4][162] 	= partial_clause_prev[4][162] & 1'b1;
			partial_clause[4][163] 	= partial_clause_prev[4][163] & 1'b1;
			partial_clause[4][164] 	= partial_clause_prev[4][164] & 1'b1;
			partial_clause[4][165] 	= partial_clause_prev[4][165] & 1'b1;
			partial_clause[4][166] 	= partial_clause_prev[4][166] & 1'b1;
			partial_clause[4][167] 	= partial_clause_prev[4][167] & 1'b1;
			partial_clause[4][168] 	= partial_clause_prev[4][168] & 1'b1;
			partial_clause[4][169] 	= partial_clause_prev[4][169] & 1'b1;
			partial_clause[4][170] 	= partial_clause_prev[4][170] & 1'b1;
			partial_clause[4][171] 	= partial_clause_prev[4][171] & 1'b1;
			partial_clause[4][172] 	= partial_clause_prev[4][172] & 1'b1;
			partial_clause[4][173] 	= partial_clause_prev[4][173] & 1'b1;
			partial_clause[4][174] 	= partial_clause_prev[4][174] & 1'b1;
			partial_clause[4][175] 	= partial_clause_prev[4][175] & 1'b1;
			partial_clause[4][176] 	= partial_clause_prev[4][176] & 1'b1;
			partial_clause[4][177] 	= partial_clause_prev[4][177] & 1'b1;
			partial_clause[4][178] 	= partial_clause_prev[4][178] & 1'b1;
			partial_clause[4][179] 	= partial_clause_prev[4][179] & 1'b1;
			partial_clause[4][180] 	= partial_clause_prev[4][180] & 1'b1;
			partial_clause[4][181] 	= partial_clause_prev[4][181] & x[53];
			partial_clause[4][182] 	= partial_clause_prev[4][182] & 1'b1;
			partial_clause[4][183] 	= partial_clause_prev[4][183] & ~x[26];
			partial_clause[4][184] 	= partial_clause_prev[4][184] & 1'b1;
			partial_clause[4][185] 	= partial_clause_prev[4][185] & 1'b1;
			partial_clause[4][186] 	= partial_clause_prev[4][186] & 1'b1;
			partial_clause[4][187] 	= partial_clause_prev[4][187] & 1'b1;
			partial_clause[4][188] 	= partial_clause_prev[4][188] & 1'b1;
			partial_clause[4][189] 	= partial_clause_prev[4][189] & 1'b1;
			partial_clause[4][190] 	= partial_clause_prev[4][190] & 1'b1;
			partial_clause[4][191] 	= partial_clause_prev[4][191] & 1'b1;
			partial_clause[4][192] 	= partial_clause_prev[4][192] & 1'b1;
			partial_clause[4][193] 	= partial_clause_prev[4][193] & 1'b1;
			partial_clause[4][194] 	= partial_clause_prev[4][194] & ~x[32];
			partial_clause[4][195] 	= partial_clause_prev[4][195] & 1'b1;
			partial_clause[4][196] 	= partial_clause_prev[4][196] & 1'b1;
			partial_clause[4][197] 	= partial_clause_prev[4][197] & 1'b1;
			partial_clause[4][198] 	= partial_clause_prev[4][198] & 1'b1;
			partial_clause[4][199] 	= partial_clause_prev[4][199] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & ~x[56];
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & x[57];
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & x[6];
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & ~x[56];
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & ~x[21];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & x[34];
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & x[63];
			partial_clause[5][38] 	= partial_clause_prev[5][38] & x[6];
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & x[29];
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & ~x[53] & ~x[56];
			partial_clause[5][47] 	= partial_clause_prev[5][47] & x[35];
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & ~x[30];
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & ~x[0];
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & ~x[0];
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & x[32];
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & ~x[3] & ~x[27] & ~x[55] & ~x[56];
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & ~x[30] & ~x[31];
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & x[9];
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & x[60];
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & x[33];
			partial_clause[5][98] 	= partial_clause_prev[5][98] & x[57];
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			partial_clause[5][100] 	= partial_clause_prev[5][100] & 1'b1;
			partial_clause[5][101] 	= partial_clause_prev[5][101] & 1'b1;
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & 1'b1;
			partial_clause[5][104] 	= partial_clause_prev[5][104] & 1'b1;
			partial_clause[5][105] 	= partial_clause_prev[5][105] & 1'b1;
			partial_clause[5][106] 	= partial_clause_prev[5][106] & 1'b1;
			partial_clause[5][107] 	= partial_clause_prev[5][107] & 1'b1;
			partial_clause[5][108] 	= partial_clause_prev[5][108] & 1'b1;
			partial_clause[5][109] 	= partial_clause_prev[5][109] & 1'b1;
			partial_clause[5][110] 	= partial_clause_prev[5][110] & 1'b1;
			partial_clause[5][111] 	= partial_clause_prev[5][111] & 1'b1;
			partial_clause[5][112] 	= partial_clause_prev[5][112] & 1'b1;
			partial_clause[5][113] 	= partial_clause_prev[5][113] & 1'b1;
			partial_clause[5][114] 	= partial_clause_prev[5][114] & 1'b1;
			partial_clause[5][115] 	= partial_clause_prev[5][115] & 1'b1;
			partial_clause[5][116] 	= partial_clause_prev[5][116] & 1'b1;
			partial_clause[5][117] 	= partial_clause_prev[5][117] & 1'b1;
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & 1'b1;
			partial_clause[5][120] 	= partial_clause_prev[5][120] & 1'b1;
			partial_clause[5][121] 	= partial_clause_prev[5][121] & 1'b1;
			partial_clause[5][122] 	= partial_clause_prev[5][122] & 1'b1;
			partial_clause[5][123] 	= partial_clause_prev[5][123] & 1'b1;
			partial_clause[5][124] 	= partial_clause_prev[5][124] & 1'b1;
			partial_clause[5][125] 	= partial_clause_prev[5][125] & 1'b1;
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & 1'b1;
			partial_clause[5][128] 	= partial_clause_prev[5][128] & 1'b1;
			partial_clause[5][129] 	= partial_clause_prev[5][129] & 1'b1;
			partial_clause[5][130] 	= partial_clause_prev[5][130] & 1'b1;
			partial_clause[5][131] 	= partial_clause_prev[5][131] & 1'b1;
			partial_clause[5][132] 	= partial_clause_prev[5][132] & ~x[59];
			partial_clause[5][133] 	= partial_clause_prev[5][133] & 1'b1;
			partial_clause[5][134] 	= partial_clause_prev[5][134] & 1'b1;
			partial_clause[5][135] 	= partial_clause_prev[5][135] & 1'b1;
			partial_clause[5][136] 	= partial_clause_prev[5][136] & 1'b1;
			partial_clause[5][137] 	= partial_clause_prev[5][137] & 1'b1;
			partial_clause[5][138] 	= partial_clause_prev[5][138] & 1'b1;
			partial_clause[5][139] 	= partial_clause_prev[5][139] & 1'b1;
			partial_clause[5][140] 	= partial_clause_prev[5][140] & 1'b1;
			partial_clause[5][141] 	= partial_clause_prev[5][141] & 1'b1;
			partial_clause[5][142] 	= partial_clause_prev[5][142] & 1'b1;
			partial_clause[5][143] 	= partial_clause_prev[5][143] & 1'b1;
			partial_clause[5][144] 	= partial_clause_prev[5][144] & 1'b1;
			partial_clause[5][145] 	= partial_clause_prev[5][145] & 1'b1;
			partial_clause[5][146] 	= partial_clause_prev[5][146] & 1'b1;
			partial_clause[5][147] 	= partial_clause_prev[5][147] & 1'b1;
			partial_clause[5][148] 	= partial_clause_prev[5][148] & 1'b1;
			partial_clause[5][149] 	= partial_clause_prev[5][149] & 1'b1;
			partial_clause[5][150] 	= partial_clause_prev[5][150] & x[17];
			partial_clause[5][151] 	= partial_clause_prev[5][151] & 1'b1;
			partial_clause[5][152] 	= partial_clause_prev[5][152] & ~x[32];
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & 1'b1;
			partial_clause[5][155] 	= partial_clause_prev[5][155] & 1'b1;
			partial_clause[5][156] 	= partial_clause_prev[5][156] & 1'b1;
			partial_clause[5][157] 	= partial_clause_prev[5][157] & 1'b1;
			partial_clause[5][158] 	= partial_clause_prev[5][158] & 1'b1;
			partial_clause[5][159] 	= partial_clause_prev[5][159] & 1'b1;
			partial_clause[5][160] 	= partial_clause_prev[5][160] & 1'b1;
			partial_clause[5][161] 	= partial_clause_prev[5][161] & 1'b1;
			partial_clause[5][162] 	= partial_clause_prev[5][162] & 1'b1;
			partial_clause[5][163] 	= partial_clause_prev[5][163] & 1'b1;
			partial_clause[5][164] 	= partial_clause_prev[5][164] & 1'b1;
			partial_clause[5][165] 	= partial_clause_prev[5][165] & 1'b1;
			partial_clause[5][166] 	= partial_clause_prev[5][166] & 1'b1;
			partial_clause[5][167] 	= partial_clause_prev[5][167] & 1'b1;
			partial_clause[5][168] 	= partial_clause_prev[5][168] & 1'b1;
			partial_clause[5][169] 	= partial_clause_prev[5][169] & 1'b1;
			partial_clause[5][170] 	= partial_clause_prev[5][170] & 1'b1;
			partial_clause[5][171] 	= partial_clause_prev[5][171] & 1'b1;
			partial_clause[5][172] 	= partial_clause_prev[5][172] & 1'b1;
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & 1'b1;
			partial_clause[5][175] 	= partial_clause_prev[5][175] & 1'b1;
			partial_clause[5][176] 	= partial_clause_prev[5][176] & 1'b1;
			partial_clause[5][177] 	= partial_clause_prev[5][177] & 1'b1;
			partial_clause[5][178] 	= partial_clause_prev[5][178] & 1'b1;
			partial_clause[5][179] 	= partial_clause_prev[5][179] & ~x[32] & ~x[61];
			partial_clause[5][180] 	= partial_clause_prev[5][180] & ~x[35];
			partial_clause[5][181] 	= partial_clause_prev[5][181] & ~x[60];
			partial_clause[5][182] 	= partial_clause_prev[5][182] & 1'b1;
			partial_clause[5][183] 	= partial_clause_prev[5][183] & 1'b1;
			partial_clause[5][184] 	= partial_clause_prev[5][184] & 1'b1;
			partial_clause[5][185] 	= partial_clause_prev[5][185] & 1'b1;
			partial_clause[5][186] 	= partial_clause_prev[5][186] & 1'b1;
			partial_clause[5][187] 	= partial_clause_prev[5][187] & 1'b1;
			partial_clause[5][188] 	= partial_clause_prev[5][188] & 1'b1;
			partial_clause[5][189] 	= partial_clause_prev[5][189] & 1'b1;
			partial_clause[5][190] 	= partial_clause_prev[5][190] & ~x[63];
			partial_clause[5][191] 	= partial_clause_prev[5][191] & 1'b1;
			partial_clause[5][192] 	= partial_clause_prev[5][192] & 1'b1;
			partial_clause[5][193] 	= partial_clause_prev[5][193] & 1'b1;
			partial_clause[5][194] 	= partial_clause_prev[5][194] & 1'b1;
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & 1'b1;
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & 1'b1;
			partial_clause[5][199] 	= partial_clause_prev[5][199] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & ~x[25];
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & x[2];
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & ~x[48];
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & ~x[59];
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & ~x[28];
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & ~x[21] & ~x[24];
			partial_clause[6][20] 	= partial_clause_prev[6][20] & ~x[22] & ~x[23];
			partial_clause[6][21] 	= partial_clause_prev[6][21] & ~x[20] & ~x[49];
			partial_clause[6][22] 	= partial_clause_prev[6][22] & ~x[27];
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & ~x[25];
			partial_clause[6][37] 	= partial_clause_prev[6][37] & x[40];
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & ~x[52];
			partial_clause[6][42] 	= partial_clause_prev[6][42] & ~x[61];
			partial_clause[6][43] 	= partial_clause_prev[6][43] & x[7];
			partial_clause[6][44] 	= partial_clause_prev[6][44] & ~x[60];
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & ~x[24] & ~x[52];
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & ~x[51];
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & x[1] & ~x[25];
			partial_clause[6][56] 	= partial_clause_prev[6][56] & ~x[30] & ~x[60];
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & ~x[22];
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & ~x[58];
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & x[55];
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & ~x[24];
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & x[35];
			partial_clause[6][79] 	= partial_clause_prev[6][79] & ~x[30] & ~x[57] & ~x[61];
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & ~x[53];
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & ~x[28] & ~x[29];
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & ~x[57] & ~x[60];
			partial_clause[6][94] 	= partial_clause_prev[6][94] & x[4];
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & x[39];
			partial_clause[6][97] 	= partial_clause_prev[6][97] & ~x[58];
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			partial_clause[6][100] 	= partial_clause_prev[6][100] & 1'b1;
			partial_clause[6][101] 	= partial_clause_prev[6][101] & 1'b1;
			partial_clause[6][102] 	= partial_clause_prev[6][102] & 1'b1;
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & 1'b1;
			partial_clause[6][105] 	= partial_clause_prev[6][105] & 1'b1;
			partial_clause[6][106] 	= partial_clause_prev[6][106] & 1'b1;
			partial_clause[6][107] 	= partial_clause_prev[6][107] & 1'b1;
			partial_clause[6][108] 	= partial_clause_prev[6][108] & 1'b1;
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & 1'b1;
			partial_clause[6][111] 	= partial_clause_prev[6][111] & 1'b1;
			partial_clause[6][112] 	= partial_clause_prev[6][112] & ~x[1];
			partial_clause[6][113] 	= partial_clause_prev[6][113] & 1'b1;
			partial_clause[6][114] 	= partial_clause_prev[6][114] & 1'b1;
			partial_clause[6][115] 	= partial_clause_prev[6][115] & 1'b1;
			partial_clause[6][116] 	= partial_clause_prev[6][116] & 1'b1;
			partial_clause[6][117] 	= partial_clause_prev[6][117] & 1'b1;
			partial_clause[6][118] 	= partial_clause_prev[6][118] & ~x[3] & ~x[5] & ~x[6] & ~x[35];
			partial_clause[6][119] 	= partial_clause_prev[6][119] & 1'b1;
			partial_clause[6][120] 	= partial_clause_prev[6][120] & ~x[2] & ~x[4] & ~x[28];
			partial_clause[6][121] 	= partial_clause_prev[6][121] & x[27];
			partial_clause[6][122] 	= partial_clause_prev[6][122] & 1'b1;
			partial_clause[6][123] 	= partial_clause_prev[6][123] & 1'b1;
			partial_clause[6][124] 	= partial_clause_prev[6][124] & 1'b1;
			partial_clause[6][125] 	= partial_clause_prev[6][125] & 1'b1;
			partial_clause[6][126] 	= partial_clause_prev[6][126] & 1'b1;
			partial_clause[6][127] 	= partial_clause_prev[6][127] & 1'b1;
			partial_clause[6][128] 	= partial_clause_prev[6][128] & 1'b1;
			partial_clause[6][129] 	= partial_clause_prev[6][129] & 1'b1;
			partial_clause[6][130] 	= partial_clause_prev[6][130] & 1'b1;
			partial_clause[6][131] 	= partial_clause_prev[6][131] & 1'b1;
			partial_clause[6][132] 	= partial_clause_prev[6][132] & 1'b1;
			partial_clause[6][133] 	= partial_clause_prev[6][133] & 1'b1;
			partial_clause[6][134] 	= partial_clause_prev[6][134] & 1'b1;
			partial_clause[6][135] 	= partial_clause_prev[6][135] & 1'b1;
			partial_clause[6][136] 	= partial_clause_prev[6][136] & 1'b1;
			partial_clause[6][137] 	= partial_clause_prev[6][137] & 1'b1;
			partial_clause[6][138] 	= partial_clause_prev[6][138] & 1'b1;
			partial_clause[6][139] 	= partial_clause_prev[6][139] & ~x[3];
			partial_clause[6][140] 	= partial_clause_prev[6][140] & 1'b1;
			partial_clause[6][141] 	= partial_clause_prev[6][141] & 1'b1;
			partial_clause[6][142] 	= partial_clause_prev[6][142] & 1'b1;
			partial_clause[6][143] 	= partial_clause_prev[6][143] & 1'b1;
			partial_clause[6][144] 	= partial_clause_prev[6][144] & 1'b1;
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & 1'b1;
			partial_clause[6][147] 	= partial_clause_prev[6][147] & 1'b1;
			partial_clause[6][148] 	= partial_clause_prev[6][148] & 1'b1;
			partial_clause[6][149] 	= partial_clause_prev[6][149] & 1'b1;
			partial_clause[6][150] 	= partial_clause_prev[6][150] & 1'b1;
			partial_clause[6][151] 	= partial_clause_prev[6][151] & 1'b1;
			partial_clause[6][152] 	= partial_clause_prev[6][152] & 1'b1;
			partial_clause[6][153] 	= partial_clause_prev[6][153] & 1'b1;
			partial_clause[6][154] 	= partial_clause_prev[6][154] & 1'b1;
			partial_clause[6][155] 	= partial_clause_prev[6][155] & 1'b1;
			partial_clause[6][156] 	= partial_clause_prev[6][156] & x[56];
			partial_clause[6][157] 	= partial_clause_prev[6][157] & 1'b1;
			partial_clause[6][158] 	= partial_clause_prev[6][158] & x[27];
			partial_clause[6][159] 	= partial_clause_prev[6][159] & 1'b1;
			partial_clause[6][160] 	= partial_clause_prev[6][160] & 1'b1;
			partial_clause[6][161] 	= partial_clause_prev[6][161] & 1'b1;
			partial_clause[6][162] 	= partial_clause_prev[6][162] & 1'b1;
			partial_clause[6][163] 	= partial_clause_prev[6][163] & 1'b1;
			partial_clause[6][164] 	= partial_clause_prev[6][164] & 1'b1;
			partial_clause[6][165] 	= partial_clause_prev[6][165] & 1'b1;
			partial_clause[6][166] 	= partial_clause_prev[6][166] & 1'b1;
			partial_clause[6][167] 	= partial_clause_prev[6][167] & 1'b1;
			partial_clause[6][168] 	= partial_clause_prev[6][168] & ~x[5] & ~x[29];
			partial_clause[6][169] 	= partial_clause_prev[6][169] & 1'b1;
			partial_clause[6][170] 	= partial_clause_prev[6][170] & 1'b1;
			partial_clause[6][171] 	= partial_clause_prev[6][171] & 1'b1;
			partial_clause[6][172] 	= partial_clause_prev[6][172] & 1'b1;
			partial_clause[6][173] 	= partial_clause_prev[6][173] & 1'b1;
			partial_clause[6][174] 	= partial_clause_prev[6][174] & 1'b1;
			partial_clause[6][175] 	= partial_clause_prev[6][175] & 1'b1;
			partial_clause[6][176] 	= partial_clause_prev[6][176] & 1'b1;
			partial_clause[6][177] 	= partial_clause_prev[6][177] & 1'b1;
			partial_clause[6][178] 	= partial_clause_prev[6][178] & 1'b1;
			partial_clause[6][179] 	= partial_clause_prev[6][179] & x[57];
			partial_clause[6][180] 	= partial_clause_prev[6][180] & 1'b1;
			partial_clause[6][181] 	= partial_clause_prev[6][181] & 1'b1;
			partial_clause[6][182] 	= partial_clause_prev[6][182] & 1'b1;
			partial_clause[6][183] 	= partial_clause_prev[6][183] & 1'b1;
			partial_clause[6][184] 	= partial_clause_prev[6][184] & 1'b1;
			partial_clause[6][185] 	= partial_clause_prev[6][185] & 1'b1;
			partial_clause[6][186] 	= partial_clause_prev[6][186] & ~x[4] & ~x[33];
			partial_clause[6][187] 	= partial_clause_prev[6][187] & ~x[8] & ~x[35];
			partial_clause[6][188] 	= partial_clause_prev[6][188] & 1'b1;
			partial_clause[6][189] 	= partial_clause_prev[6][189] & 1'b1;
			partial_clause[6][190] 	= partial_clause_prev[6][190] & 1'b1;
			partial_clause[6][191] 	= partial_clause_prev[6][191] & 1'b1;
			partial_clause[6][192] 	= partial_clause_prev[6][192] & ~x[62];
			partial_clause[6][193] 	= partial_clause_prev[6][193] & 1'b1;
			partial_clause[6][194] 	= partial_clause_prev[6][194] & ~x[7];
			partial_clause[6][195] 	= partial_clause_prev[6][195] & 1'b1;
			partial_clause[6][196] 	= partial_clause_prev[6][196] & x[50];
			partial_clause[6][197] 	= partial_clause_prev[6][197] & 1'b1;
			partial_clause[6][198] 	= partial_clause_prev[6][198] & 1'b1;
			partial_clause[6][199] 	= partial_clause_prev[6][199] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & ~x[32] & ~x[53];
			partial_clause[7][1] 	= partial_clause_prev[7][1] & ~x[32];
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & ~x[56];
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & ~x[25];
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & ~x[23] & ~x[29];
			partial_clause[7][31] 	= partial_clause_prev[7][31] & ~x[33];
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & ~x[27];
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & ~x[56] & ~x[57];
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & x[15];
			partial_clause[7][83] 	= partial_clause_prev[7][83] & ~x[23];
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & ~x[53] & ~x[55];
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			partial_clause[7][100] 	= partial_clause_prev[7][100] & 1'b1;
			partial_clause[7][101] 	= partial_clause_prev[7][101] & ~x[49] & ~x[50];
			partial_clause[7][102] 	= partial_clause_prev[7][102] & 1'b1;
			partial_clause[7][103] 	= partial_clause_prev[7][103] & 1'b1;
			partial_clause[7][104] 	= partial_clause_prev[7][104] & 1'b1;
			partial_clause[7][105] 	= partial_clause_prev[7][105] & ~x[54];
			partial_clause[7][106] 	= partial_clause_prev[7][106] & 1'b1;
			partial_clause[7][107] 	= partial_clause_prev[7][107] & 1'b1;
			partial_clause[7][108] 	= partial_clause_prev[7][108] & ~x[53];
			partial_clause[7][109] 	= partial_clause_prev[7][109] & 1'b1;
			partial_clause[7][110] 	= partial_clause_prev[7][110] & x[25];
			partial_clause[7][111] 	= partial_clause_prev[7][111] & x[53];
			partial_clause[7][112] 	= partial_clause_prev[7][112] & 1'b1;
			partial_clause[7][113] 	= partial_clause_prev[7][113] & ~x[50];
			partial_clause[7][114] 	= partial_clause_prev[7][114] & 1'b1;
			partial_clause[7][115] 	= partial_clause_prev[7][115] & 1'b1;
			partial_clause[7][116] 	= partial_clause_prev[7][116] & x[30];
			partial_clause[7][117] 	= partial_clause_prev[7][117] & 1'b1;
			partial_clause[7][118] 	= partial_clause_prev[7][118] & 1'b1;
			partial_clause[7][119] 	= partial_clause_prev[7][119] & 1'b1;
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & 1'b1;
			partial_clause[7][123] 	= partial_clause_prev[7][123] & 1'b1;
			partial_clause[7][124] 	= partial_clause_prev[7][124] & 1'b1;
			partial_clause[7][125] 	= partial_clause_prev[7][125] & 1'b1;
			partial_clause[7][126] 	= partial_clause_prev[7][126] & 1'b1;
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & x[29];
			partial_clause[7][129] 	= partial_clause_prev[7][129] & 1'b1;
			partial_clause[7][130] 	= partial_clause_prev[7][130] & 1'b1;
			partial_clause[7][131] 	= partial_clause_prev[7][131] & 1'b1;
			partial_clause[7][132] 	= partial_clause_prev[7][132] & x[29];
			partial_clause[7][133] 	= partial_clause_prev[7][133] & 1'b1;
			partial_clause[7][134] 	= partial_clause_prev[7][134] & 1'b1;
			partial_clause[7][135] 	= partial_clause_prev[7][135] & 1'b1;
			partial_clause[7][136] 	= partial_clause_prev[7][136] & 1'b1;
			partial_clause[7][137] 	= partial_clause_prev[7][137] & ~x[51];
			partial_clause[7][138] 	= partial_clause_prev[7][138] & 1'b1;
			partial_clause[7][139] 	= partial_clause_prev[7][139] & 1'b1;
			partial_clause[7][140] 	= partial_clause_prev[7][140] & 1'b1;
			partial_clause[7][141] 	= partial_clause_prev[7][141] & 1'b1;
			partial_clause[7][142] 	= partial_clause_prev[7][142] & 1'b1;
			partial_clause[7][143] 	= partial_clause_prev[7][143] & 1'b1;
			partial_clause[7][144] 	= partial_clause_prev[7][144] & x[27];
			partial_clause[7][145] 	= partial_clause_prev[7][145] & 1'b1;
			partial_clause[7][146] 	= partial_clause_prev[7][146] & 1'b1;
			partial_clause[7][147] 	= partial_clause_prev[7][147] & 1'b1;
			partial_clause[7][148] 	= partial_clause_prev[7][148] & x[27];
			partial_clause[7][149] 	= partial_clause_prev[7][149] & x[30];
			partial_clause[7][150] 	= partial_clause_prev[7][150] & 1'b1;
			partial_clause[7][151] 	= partial_clause_prev[7][151] & 1'b1;
			partial_clause[7][152] 	= partial_clause_prev[7][152] & 1'b1;
			partial_clause[7][153] 	= partial_clause_prev[7][153] & 1'b1;
			partial_clause[7][154] 	= partial_clause_prev[7][154] & 1'b1;
			partial_clause[7][155] 	= partial_clause_prev[7][155] & 1'b1;
			partial_clause[7][156] 	= partial_clause_prev[7][156] & x[25];
			partial_clause[7][157] 	= partial_clause_prev[7][157] & 1'b1;
			partial_clause[7][158] 	= partial_clause_prev[7][158] & 1'b1;
			partial_clause[7][159] 	= partial_clause_prev[7][159] & 1'b1;
			partial_clause[7][160] 	= partial_clause_prev[7][160] & 1'b1;
			partial_clause[7][161] 	= partial_clause_prev[7][161] & x[53];
			partial_clause[7][162] 	= partial_clause_prev[7][162] & 1'b1;
			partial_clause[7][163] 	= partial_clause_prev[7][163] & 1'b1;
			partial_clause[7][164] 	= partial_clause_prev[7][164] & 1'b1;
			partial_clause[7][165] 	= partial_clause_prev[7][165] & x[31];
			partial_clause[7][166] 	= partial_clause_prev[7][166] & 1'b1;
			partial_clause[7][167] 	= partial_clause_prev[7][167] & 1'b1;
			partial_clause[7][168] 	= partial_clause_prev[7][168] & 1'b1;
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & 1'b1;
			partial_clause[7][171] 	= partial_clause_prev[7][171] & 1'b1;
			partial_clause[7][172] 	= partial_clause_prev[7][172] & 1'b1;
			partial_clause[7][173] 	= partial_clause_prev[7][173] & 1'b1;
			partial_clause[7][174] 	= partial_clause_prev[7][174] & x[28];
			partial_clause[7][175] 	= partial_clause_prev[7][175] & 1'b1;
			partial_clause[7][176] 	= partial_clause_prev[7][176] & x[31];
			partial_clause[7][177] 	= partial_clause_prev[7][177] & 1'b1;
			partial_clause[7][178] 	= partial_clause_prev[7][178] & 1'b1;
			partial_clause[7][179] 	= partial_clause_prev[7][179] & 1'b1;
			partial_clause[7][180] 	= partial_clause_prev[7][180] & 1'b1;
			partial_clause[7][181] 	= partial_clause_prev[7][181] & 1'b1;
			partial_clause[7][182] 	= partial_clause_prev[7][182] & 1'b1;
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & 1'b1;
			partial_clause[7][185] 	= partial_clause_prev[7][185] & 1'b1;
			partial_clause[7][186] 	= partial_clause_prev[7][186] & 1'b1;
			partial_clause[7][187] 	= partial_clause_prev[7][187] & 1'b1;
			partial_clause[7][188] 	= partial_clause_prev[7][188] & 1'b1;
			partial_clause[7][189] 	= partial_clause_prev[7][189] & 1'b1;
			partial_clause[7][190] 	= partial_clause_prev[7][190] & 1'b1;
			partial_clause[7][191] 	= partial_clause_prev[7][191] & 1'b1;
			partial_clause[7][192] 	= partial_clause_prev[7][192] & 1'b1;
			partial_clause[7][193] 	= partial_clause_prev[7][193] & 1'b1;
			partial_clause[7][194] 	= partial_clause_prev[7][194] & x[34];
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & 1'b1;
			partial_clause[7][197] 	= partial_clause_prev[7][197] & 1'b1;
			partial_clause[7][198] 	= partial_clause_prev[7][198] & 1'b1;
			partial_clause[7][199] 	= partial_clause_prev[7][199] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & x[53];
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & ~x[32];
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & x[26];
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & ~x[47];
			partial_clause[8][17] 	= partial_clause_prev[8][17] & x[27];
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & ~x[0];
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & x[13];
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & x[14];
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & x[13];
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & x[11];
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & ~x[22];
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & ~x[49];
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & x[8];
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & x[42];
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			partial_clause[8][100] 	= partial_clause_prev[8][100] & 1'b1;
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & ~x[16] & ~x[52];
			partial_clause[8][103] 	= partial_clause_prev[8][103] & 1'b1;
			partial_clause[8][104] 	= partial_clause_prev[8][104] & 1'b1;
			partial_clause[8][105] 	= partial_clause_prev[8][105] & 1'b1;
			partial_clause[8][106] 	= partial_clause_prev[8][106] & 1'b1;
			partial_clause[8][107] 	= partial_clause_prev[8][107] & 1'b1;
			partial_clause[8][108] 	= partial_clause_prev[8][108] & 1'b1;
			partial_clause[8][109] 	= partial_clause_prev[8][109] & 1'b1;
			partial_clause[8][110] 	= partial_clause_prev[8][110] & 1'b1;
			partial_clause[8][111] 	= partial_clause_prev[8][111] & 1'b1;
			partial_clause[8][112] 	= partial_clause_prev[8][112] & 1'b1;
			partial_clause[8][113] 	= partial_clause_prev[8][113] & 1'b1;
			partial_clause[8][114] 	= partial_clause_prev[8][114] & ~x[0] & ~x[27] & ~x[55] & ~x[56];
			partial_clause[8][115] 	= partial_clause_prev[8][115] & x[46];
			partial_clause[8][116] 	= partial_clause_prev[8][116] & 1'b1;
			partial_clause[8][117] 	= partial_clause_prev[8][117] & 1'b1;
			partial_clause[8][118] 	= partial_clause_prev[8][118] & 1'b1;
			partial_clause[8][119] 	= partial_clause_prev[8][119] & 1'b1;
			partial_clause[8][120] 	= partial_clause_prev[8][120] & 1'b1;
			partial_clause[8][121] 	= partial_clause_prev[8][121] & 1'b1;
			partial_clause[8][122] 	= partial_clause_prev[8][122] & 1'b1;
			partial_clause[8][123] 	= partial_clause_prev[8][123] & 1'b1;
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & 1'b1;
			partial_clause[8][126] 	= partial_clause_prev[8][126] & 1'b1;
			partial_clause[8][127] 	= partial_clause_prev[8][127] & 1'b1;
			partial_clause[8][128] 	= partial_clause_prev[8][128] & 1'b1;
			partial_clause[8][129] 	= partial_clause_prev[8][129] & 1'b1;
			partial_clause[8][130] 	= partial_clause_prev[8][130] & 1'b1;
			partial_clause[8][131] 	= partial_clause_prev[8][131] & 1'b1;
			partial_clause[8][132] 	= partial_clause_prev[8][132] & ~x[29] & ~x[52];
			partial_clause[8][133] 	= partial_clause_prev[8][133] & 1'b1;
			partial_clause[8][134] 	= partial_clause_prev[8][134] & x[20];
			partial_clause[8][135] 	= partial_clause_prev[8][135] & 1'b1;
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & 1'b1;
			partial_clause[8][138] 	= partial_clause_prev[8][138] & 1'b1;
			partial_clause[8][139] 	= partial_clause_prev[8][139] & ~x[30];
			partial_clause[8][140] 	= partial_clause_prev[8][140] & 1'b1;
			partial_clause[8][141] 	= partial_clause_prev[8][141] & 1'b1;
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & 1'b1;
			partial_clause[8][144] 	= partial_clause_prev[8][144] & 1'b1;
			partial_clause[8][145] 	= partial_clause_prev[8][145] & 1'b1;
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & 1'b1;
			partial_clause[8][148] 	= partial_clause_prev[8][148] & 1'b1;
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & 1'b1;
			partial_clause[8][151] 	= partial_clause_prev[8][151] & 1'b1;
			partial_clause[8][152] 	= partial_clause_prev[8][152] & 1'b1;
			partial_clause[8][153] 	= partial_clause_prev[8][153] & 1'b1;
			partial_clause[8][154] 	= partial_clause_prev[8][154] & 1'b1;
			partial_clause[8][155] 	= partial_clause_prev[8][155] & 1'b1;
			partial_clause[8][156] 	= partial_clause_prev[8][156] & 1'b1;
			partial_clause[8][157] 	= partial_clause_prev[8][157] & 1'b1;
			partial_clause[8][158] 	= partial_clause_prev[8][158] & 1'b1;
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & x[20];
			partial_clause[8][161] 	= partial_clause_prev[8][161] & 1'b1;
			partial_clause[8][162] 	= partial_clause_prev[8][162] & 1'b1;
			partial_clause[8][163] 	= partial_clause_prev[8][163] & 1'b1;
			partial_clause[8][164] 	= partial_clause_prev[8][164] & 1'b1;
			partial_clause[8][165] 	= partial_clause_prev[8][165] & 1'b1;
			partial_clause[8][166] 	= partial_clause_prev[8][166] & 1'b1;
			partial_clause[8][167] 	= partial_clause_prev[8][167] & 1'b1;
			partial_clause[8][168] 	= partial_clause_prev[8][168] & 1'b1;
			partial_clause[8][169] 	= partial_clause_prev[8][169] & 1'b1;
			partial_clause[8][170] 	= partial_clause_prev[8][170] & 1'b1;
			partial_clause[8][171] 	= partial_clause_prev[8][171] & 1'b1;
			partial_clause[8][172] 	= partial_clause_prev[8][172] & 1'b1;
			partial_clause[8][173] 	= partial_clause_prev[8][173] & 1'b1;
			partial_clause[8][174] 	= partial_clause_prev[8][174] & 1'b1;
			partial_clause[8][175] 	= partial_clause_prev[8][175] & 1'b1;
			partial_clause[8][176] 	= partial_clause_prev[8][176] & x[18];
			partial_clause[8][177] 	= partial_clause_prev[8][177] & 1'b1;
			partial_clause[8][178] 	= partial_clause_prev[8][178] & x[47];
			partial_clause[8][179] 	= partial_clause_prev[8][179] & 1'b1;
			partial_clause[8][180] 	= partial_clause_prev[8][180] & 1'b1;
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & 1'b1;
			partial_clause[8][183] 	= partial_clause_prev[8][183] & 1'b1;
			partial_clause[8][184] 	= partial_clause_prev[8][184] & 1'b1;
			partial_clause[8][185] 	= partial_clause_prev[8][185] & 1'b1;
			partial_clause[8][186] 	= partial_clause_prev[8][186] & 1'b1;
			partial_clause[8][187] 	= partial_clause_prev[8][187] & 1'b1;
			partial_clause[8][188] 	= partial_clause_prev[8][188] & 1'b1;
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & 1'b1;
			partial_clause[8][191] 	= partial_clause_prev[8][191] & 1'b1;
			partial_clause[8][192] 	= partial_clause_prev[8][192] & 1'b1;
			partial_clause[8][193] 	= partial_clause_prev[8][193] & 1'b1;
			partial_clause[8][194] 	= partial_clause_prev[8][194] & ~x[52];
			partial_clause[8][195] 	= partial_clause_prev[8][195] & 1'b1;
			partial_clause[8][196] 	= partial_clause_prev[8][196] & 1'b1;
			partial_clause[8][197] 	= partial_clause_prev[8][197] & 1'b1;
			partial_clause[8][198] 	= partial_clause_prev[8][198] & 1'b1;
			partial_clause[8][199] 	= partial_clause_prev[8][199] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & ~x[26] & ~x[28];
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & x[54];
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & x[56];
			partial_clause[9][35] 	= partial_clause_prev[9][35] & ~x[62];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & ~x[24] & ~x[50];
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & ~x[50] & ~x[59];
			partial_clause[9][49] 	= partial_clause_prev[9][49] & ~x[27];
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & ~x[27] & ~x[28];
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & ~x[26];
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & ~x[26];
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & ~x[26];
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & ~x[27] & ~x[28];
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & ~x[3] & ~x[63];
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & x[12];
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & ~x[26];
			partial_clause[9][100] 	= partial_clause_prev[9][100] & 1'b1;
			partial_clause[9][101] 	= partial_clause_prev[9][101] & ~x[56];
			partial_clause[9][102] 	= partial_clause_prev[9][102] & x[27];
			partial_clause[9][103] 	= partial_clause_prev[9][103] & x[62];
			partial_clause[9][104] 	= partial_clause_prev[9][104] & x[49];
			partial_clause[9][105] 	= partial_clause_prev[9][105] & 1'b1;
			partial_clause[9][106] 	= partial_clause_prev[9][106] & x[62];
			partial_clause[9][107] 	= partial_clause_prev[9][107] & x[29];
			partial_clause[9][108] 	= partial_clause_prev[9][108] & 1'b1;
			partial_clause[9][109] 	= partial_clause_prev[9][109] & ~x[55];
			partial_clause[9][110] 	= partial_clause_prev[9][110] & 1'b1;
			partial_clause[9][111] 	= partial_clause_prev[9][111] & 1'b1;
			partial_clause[9][112] 	= partial_clause_prev[9][112] & x[0];
			partial_clause[9][113] 	= partial_clause_prev[9][113] & 1'b1;
			partial_clause[9][114] 	= partial_clause_prev[9][114] & 1'b1;
			partial_clause[9][115] 	= partial_clause_prev[9][115] & 1'b1;
			partial_clause[9][116] 	= partial_clause_prev[9][116] & 1'b1;
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & ~x[56];
			partial_clause[9][119] 	= partial_clause_prev[9][119] & 1'b1;
			partial_clause[9][120] 	= partial_clause_prev[9][120] & x[30];
			partial_clause[9][121] 	= partial_clause_prev[9][121] & x[1];
			partial_clause[9][122] 	= partial_clause_prev[9][122] & 1'b1;
			partial_clause[9][123] 	= partial_clause_prev[9][123] & x[32];
			partial_clause[9][124] 	= partial_clause_prev[9][124] & 1'b1;
			partial_clause[9][125] 	= partial_clause_prev[9][125] & 1'b1;
			partial_clause[9][126] 	= partial_clause_prev[9][126] & 1'b1;
			partial_clause[9][127] 	= partial_clause_prev[9][127] & 1'b1;
			partial_clause[9][128] 	= partial_clause_prev[9][128] & 1'b1;
			partial_clause[9][129] 	= partial_clause_prev[9][129] & 1'b1;
			partial_clause[9][130] 	= partial_clause_prev[9][130] & 1'b1;
			partial_clause[9][131] 	= partial_clause_prev[9][131] & 1'b1;
			partial_clause[9][132] 	= partial_clause_prev[9][132] & 1'b1;
			partial_clause[9][133] 	= partial_clause_prev[9][133] & 1'b1;
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & x[30];
			partial_clause[9][138] 	= partial_clause_prev[9][138] & x[29];
			partial_clause[9][139] 	= partial_clause_prev[9][139] & 1'b1;
			partial_clause[9][140] 	= partial_clause_prev[9][140] & 1'b1;
			partial_clause[9][141] 	= partial_clause_prev[9][141] & 1'b1;
			partial_clause[9][142] 	= partial_clause_prev[9][142] & 1'b1;
			partial_clause[9][143] 	= partial_clause_prev[9][143] & 1'b1;
			partial_clause[9][144] 	= partial_clause_prev[9][144] & ~x[57];
			partial_clause[9][145] 	= partial_clause_prev[9][145] & x[31];
			partial_clause[9][146] 	= partial_clause_prev[9][146] & x[21];
			partial_clause[9][147] 	= partial_clause_prev[9][147] & 1'b1;
			partial_clause[9][148] 	= partial_clause_prev[9][148] & 1'b1;
			partial_clause[9][149] 	= partial_clause_prev[9][149] & 1'b1;
			partial_clause[9][150] 	= partial_clause_prev[9][150] & 1'b1;
			partial_clause[9][151] 	= partial_clause_prev[9][151] & 1'b1;
			partial_clause[9][152] 	= partial_clause_prev[9][152] & x[2];
			partial_clause[9][153] 	= partial_clause_prev[9][153] & 1'b1;
			partial_clause[9][154] 	= partial_clause_prev[9][154] & 1'b1;
			partial_clause[9][155] 	= partial_clause_prev[9][155] & ~x[55];
			partial_clause[9][156] 	= partial_clause_prev[9][156] & 1'b1;
			partial_clause[9][157] 	= partial_clause_prev[9][157] & 1'b1;
			partial_clause[9][158] 	= partial_clause_prev[9][158] & 1'b1;
			partial_clause[9][159] 	= partial_clause_prev[9][159] & 1'b1;
			partial_clause[9][160] 	= partial_clause_prev[9][160] & 1'b1;
			partial_clause[9][161] 	= partial_clause_prev[9][161] & 1'b1;
			partial_clause[9][162] 	= partial_clause_prev[9][162] & 1'b1;
			partial_clause[9][163] 	= partial_clause_prev[9][163] & x[3];
			partial_clause[9][164] 	= partial_clause_prev[9][164] & ~x[55];
			partial_clause[9][165] 	= partial_clause_prev[9][165] & 1'b1;
			partial_clause[9][166] 	= partial_clause_prev[9][166] & 1'b1;
			partial_clause[9][167] 	= partial_clause_prev[9][167] & 1'b1;
			partial_clause[9][168] 	= partial_clause_prev[9][168] & 1'b1;
			partial_clause[9][169] 	= partial_clause_prev[9][169] & 1'b1;
			partial_clause[9][170] 	= partial_clause_prev[9][170] & 1'b1;
			partial_clause[9][171] 	= partial_clause_prev[9][171] & 1'b1;
			partial_clause[9][172] 	= partial_clause_prev[9][172] & 1'b1;
			partial_clause[9][173] 	= partial_clause_prev[9][173] & 1'b1;
			partial_clause[9][174] 	= partial_clause_prev[9][174] & x[31];
			partial_clause[9][175] 	= partial_clause_prev[9][175] & ~x[27] & ~x[55];
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & 1'b1;
			partial_clause[9][178] 	= partial_clause_prev[9][178] & x[22];
			partial_clause[9][179] 	= partial_clause_prev[9][179] & 1'b1;
			partial_clause[9][180] 	= partial_clause_prev[9][180] & 1'b1;
			partial_clause[9][181] 	= partial_clause_prev[9][181] & 1'b1;
			partial_clause[9][182] 	= partial_clause_prev[9][182] & 1'b1;
			partial_clause[9][183] 	= partial_clause_prev[9][183] & x[32];
			partial_clause[9][184] 	= partial_clause_prev[9][184] & ~x[53];
			partial_clause[9][185] 	= partial_clause_prev[9][185] & x[63];
			partial_clause[9][186] 	= partial_clause_prev[9][186] & 1'b1;
			partial_clause[9][187] 	= partial_clause_prev[9][187] & ~x[26] & ~x[54];
			partial_clause[9][188] 	= partial_clause_prev[9][188] & 1'b1;
			partial_clause[9][189] 	= partial_clause_prev[9][189] & 1'b1;
			partial_clause[9][190] 	= partial_clause_prev[9][190] & x[33];
			partial_clause[9][191] 	= partial_clause_prev[9][191] & x[21];
			partial_clause[9][192] 	= partial_clause_prev[9][192] & 1'b1;
			partial_clause[9][193] 	= partial_clause_prev[9][193] & x[48];
			partial_clause[9][194] 	= partial_clause_prev[9][194] & 1'b1;
			partial_clause[9][195] 	= partial_clause_prev[9][195] & ~x[57];
			partial_clause[9][196] 	= partial_clause_prev[9][196] & 1'b1;
			partial_clause[9][197] 	= partial_clause_prev[9][197] & x[29];
			partial_clause[9][198] 	= partial_clause_prev[9][198] & 1'b1;
			partial_clause[9][199] 	= partial_clause_prev[9][199] & 1'b1;
		end
	end
endmodule


module HCB_3 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & x[3];
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & ~x[15] & x[50];
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & x[20];
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & x[25];
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & x[24];
			partial_clause[0][28] 	= partial_clause_prev[0][28] & ~x[29];
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & x[24];
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & x[22];
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & ~x[54];
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & x[21];
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & ~x[10];
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & x[48];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & x[27];
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & x[50];
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			partial_clause[0][100] 	= partial_clause_prev[0][100] & x[37];
			partial_clause[0][101] 	= partial_clause_prev[0][101] & 1'b1;
			partial_clause[0][102] 	= partial_clause_prev[0][102] & 1'b1;
			partial_clause[0][103] 	= partial_clause_prev[0][103] & 1'b1;
			partial_clause[0][104] 	= partial_clause_prev[0][104] & 1'b1;
			partial_clause[0][105] 	= partial_clause_prev[0][105] & 1'b1;
			partial_clause[0][106] 	= partial_clause_prev[0][106] & 1'b1;
			partial_clause[0][107] 	= partial_clause_prev[0][107] & 1'b1;
			partial_clause[0][108] 	= partial_clause_prev[0][108] & 1'b1;
			partial_clause[0][109] 	= partial_clause_prev[0][109] & 1'b1;
			partial_clause[0][110] 	= partial_clause_prev[0][110] & ~x[47];
			partial_clause[0][111] 	= partial_clause_prev[0][111] & 1'b1;
			partial_clause[0][112] 	= partial_clause_prev[0][112] & 1'b1;
			partial_clause[0][113] 	= partial_clause_prev[0][113] & 1'b1;
			partial_clause[0][114] 	= partial_clause_prev[0][114] & 1'b1;
			partial_clause[0][115] 	= partial_clause_prev[0][115] & 1'b1;
			partial_clause[0][116] 	= partial_clause_prev[0][116] & 1'b1;
			partial_clause[0][117] 	= partial_clause_prev[0][117] & ~x[20] & ~x[21] & ~x[22];
			partial_clause[0][118] 	= partial_clause_prev[0][118] & 1'b1;
			partial_clause[0][119] 	= partial_clause_prev[0][119] & 1'b1;
			partial_clause[0][120] 	= partial_clause_prev[0][120] & 1'b1;
			partial_clause[0][121] 	= partial_clause_prev[0][121] & 1'b1;
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & 1'b1;
			partial_clause[0][124] 	= partial_clause_prev[0][124] & 1'b1;
			partial_clause[0][125] 	= partial_clause_prev[0][125] & 1'b1;
			partial_clause[0][126] 	= partial_clause_prev[0][126] & 1'b1;
			partial_clause[0][127] 	= partial_clause_prev[0][127] & 1'b1;
			partial_clause[0][128] 	= partial_clause_prev[0][128] & 1'b1;
			partial_clause[0][129] 	= partial_clause_prev[0][129] & 1'b1;
			partial_clause[0][130] 	= partial_clause_prev[0][130] & 1'b1;
			partial_clause[0][131] 	= partial_clause_prev[0][131] & 1'b1;
			partial_clause[0][132] 	= partial_clause_prev[0][132] & 1'b1;
			partial_clause[0][133] 	= partial_clause_prev[0][133] & 1'b1;
			partial_clause[0][134] 	= partial_clause_prev[0][134] & 1'b1;
			partial_clause[0][135] 	= partial_clause_prev[0][135] & 1'b1;
			partial_clause[0][136] 	= partial_clause_prev[0][136] & ~x[31];
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & 1'b1;
			partial_clause[0][139] 	= partial_clause_prev[0][139] & 1'b1;
			partial_clause[0][140] 	= partial_clause_prev[0][140] & 1'b1;
			partial_clause[0][141] 	= partial_clause_prev[0][141] & 1'b1;
			partial_clause[0][142] 	= partial_clause_prev[0][142] & 1'b1;
			partial_clause[0][143] 	= partial_clause_prev[0][143] & 1'b1;
			partial_clause[0][144] 	= partial_clause_prev[0][144] & 1'b1;
			partial_clause[0][145] 	= partial_clause_prev[0][145] & 1'b1;
			partial_clause[0][146] 	= partial_clause_prev[0][146] & 1'b1;
			partial_clause[0][147] 	= partial_clause_prev[0][147] & ~x[26];
			partial_clause[0][148] 	= partial_clause_prev[0][148] & x[59];
			partial_clause[0][149] 	= partial_clause_prev[0][149] & ~x[48];
			partial_clause[0][150] 	= partial_clause_prev[0][150] & 1'b1;
			partial_clause[0][151] 	= partial_clause_prev[0][151] & 1'b1;
			partial_clause[0][152] 	= partial_clause_prev[0][152] & ~x[25] & ~x[49] & ~x[51];
			partial_clause[0][153] 	= partial_clause_prev[0][153] & 1'b1;
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & 1'b1;
			partial_clause[0][156] 	= partial_clause_prev[0][156] & 1'b1;
			partial_clause[0][157] 	= partial_clause_prev[0][157] & 1'b1;
			partial_clause[0][158] 	= partial_clause_prev[0][158] & 1'b1;
			partial_clause[0][159] 	= partial_clause_prev[0][159] & 1'b1;
			partial_clause[0][160] 	= partial_clause_prev[0][160] & 1'b1;
			partial_clause[0][161] 	= partial_clause_prev[0][161] & ~x[48];
			partial_clause[0][162] 	= partial_clause_prev[0][162] & 1'b1;
			partial_clause[0][163] 	= partial_clause_prev[0][163] & 1'b1;
			partial_clause[0][164] 	= partial_clause_prev[0][164] & 1'b1;
			partial_clause[0][165] 	= partial_clause_prev[0][165] & 1'b1;
			partial_clause[0][166] 	= partial_clause_prev[0][166] & 1'b1;
			partial_clause[0][167] 	= partial_clause_prev[0][167] & 1'b1;
			partial_clause[0][168] 	= partial_clause_prev[0][168] & 1'b1;
			partial_clause[0][169] 	= partial_clause_prev[0][169] & 1'b1;
			partial_clause[0][170] 	= partial_clause_prev[0][170] & 1'b1;
			partial_clause[0][171] 	= partial_clause_prev[0][171] & x[57];
			partial_clause[0][172] 	= partial_clause_prev[0][172] & 1'b1;
			partial_clause[0][173] 	= partial_clause_prev[0][173] & ~x[54];
			partial_clause[0][174] 	= partial_clause_prev[0][174] & 1'b1;
			partial_clause[0][175] 	= partial_clause_prev[0][175] & 1'b1;
			partial_clause[0][176] 	= partial_clause_prev[0][176] & 1'b1;
			partial_clause[0][177] 	= partial_clause_prev[0][177] & 1'b1;
			partial_clause[0][178] 	= partial_clause_prev[0][178] & 1'b1;
			partial_clause[0][179] 	= partial_clause_prev[0][179] & 1'b1;
			partial_clause[0][180] 	= partial_clause_prev[0][180] & 1'b1;
			partial_clause[0][181] 	= partial_clause_prev[0][181] & 1'b1;
			partial_clause[0][182] 	= partial_clause_prev[0][182] & 1'b1;
			partial_clause[0][183] 	= partial_clause_prev[0][183] & 1'b1;
			partial_clause[0][184] 	= partial_clause_prev[0][184] & 1'b1;
			partial_clause[0][185] 	= partial_clause_prev[0][185] & 1'b1;
			partial_clause[0][186] 	= partial_clause_prev[0][186] & 1'b1;
			partial_clause[0][187] 	= partial_clause_prev[0][187] & 1'b1;
			partial_clause[0][188] 	= partial_clause_prev[0][188] & 1'b1;
			partial_clause[0][189] 	= partial_clause_prev[0][189] & 1'b1;
			partial_clause[0][190] 	= partial_clause_prev[0][190] & 1'b1;
			partial_clause[0][191] 	= partial_clause_prev[0][191] & 1'b1;
			partial_clause[0][192] 	= partial_clause_prev[0][192] & 1'b1;
			partial_clause[0][193] 	= partial_clause_prev[0][193] & 1'b1;
			partial_clause[0][194] 	= partial_clause_prev[0][194] & 1'b1;
			partial_clause[0][195] 	= partial_clause_prev[0][195] & x[11];
			partial_clause[0][196] 	= partial_clause_prev[0][196] & 1'b1;
			partial_clause[0][197] 	= partial_clause_prev[0][197] & 1'b1;
			partial_clause[0][198] 	= partial_clause_prev[0][198] & 1'b1;
			partial_clause[0][199] 	= partial_clause_prev[0][199] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[45];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & x[62];
			partial_clause[1][5] 	= partial_clause_prev[1][5] & ~x[45];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & ~x[22];
			partial_clause[1][9] 	= partial_clause_prev[1][9] & ~x[17] & ~x[45];
			partial_clause[1][10] 	= partial_clause_prev[1][10] & ~x[49];
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & ~x[23] & ~x[50];
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & ~x[23] & ~x[49];
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & ~x[12] & ~x[41];
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & x[1];
			partial_clause[1][27] 	= partial_clause_prev[1][27] & ~x[22];
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & ~x[51];
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & ~x[44] & ~x[45];
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & x[61];
			partial_clause[1][52] 	= partial_clause_prev[1][52] & ~x[17];
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & x[58];
			partial_clause[1][58] 	= partial_clause_prev[1][58] & 1'b1;
			partial_clause[1][59] 	= partial_clause_prev[1][59] & ~x[52];
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & x[3];
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & ~x[15];
			partial_clause[1][67] 	= partial_clause_prev[1][67] & x[59];
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & ~x[44];
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & ~x[25];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & ~x[19];
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & x[45] & ~x[50];
			partial_clause[1][90] 	= partial_clause_prev[1][90] & ~x[17] & ~x[45];
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & ~x[15] & ~x[45];
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			partial_clause[1][100] 	= partial_clause_prev[1][100] & 1'b1;
			partial_clause[1][101] 	= partial_clause_prev[1][101] & 1'b1;
			partial_clause[1][102] 	= partial_clause_prev[1][102] & 1'b1;
			partial_clause[1][103] 	= partial_clause_prev[1][103] & 1'b1;
			partial_clause[1][104] 	= partial_clause_prev[1][104] & 1'b1;
			partial_clause[1][105] 	= partial_clause_prev[1][105] & 1'b1;
			partial_clause[1][106] 	= partial_clause_prev[1][106] & x[15];
			partial_clause[1][107] 	= partial_clause_prev[1][107] & 1'b1;
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & 1'b1;
			partial_clause[1][110] 	= partial_clause_prev[1][110] & x[44];
			partial_clause[1][111] 	= partial_clause_prev[1][111] & 1'b1;
			partial_clause[1][112] 	= partial_clause_prev[1][112] & 1'b1;
			partial_clause[1][113] 	= partial_clause_prev[1][113] & 1'b1;
			partial_clause[1][114] 	= partial_clause_prev[1][114] & 1'b1;
			partial_clause[1][115] 	= partial_clause_prev[1][115] & 1'b1;
			partial_clause[1][116] 	= partial_clause_prev[1][116] & 1'b1;
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & x[19];
			partial_clause[1][119] 	= partial_clause_prev[1][119] & 1'b1;
			partial_clause[1][120] 	= partial_clause_prev[1][120] & x[44];
			partial_clause[1][121] 	= partial_clause_prev[1][121] & 1'b1;
			partial_clause[1][122] 	= partial_clause_prev[1][122] & 1'b1;
			partial_clause[1][123] 	= partial_clause_prev[1][123] & 1'b1;
			partial_clause[1][124] 	= partial_clause_prev[1][124] & 1'b1;
			partial_clause[1][125] 	= partial_clause_prev[1][125] & 1'b1;
			partial_clause[1][126] 	= partial_clause_prev[1][126] & 1'b1;
			partial_clause[1][127] 	= partial_clause_prev[1][127] & 1'b1;
			partial_clause[1][128] 	= partial_clause_prev[1][128] & 1'b1;
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & 1'b1;
			partial_clause[1][131] 	= partial_clause_prev[1][131] & 1'b1;
			partial_clause[1][132] 	= partial_clause_prev[1][132] & 1'b1;
			partial_clause[1][133] 	= partial_clause_prev[1][133] & 1'b1;
			partial_clause[1][134] 	= partial_clause_prev[1][134] & 1'b1;
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & 1'b1;
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & 1'b1;
			partial_clause[1][139] 	= partial_clause_prev[1][139] & 1'b1;
			partial_clause[1][140] 	= partial_clause_prev[1][140] & 1'b1;
			partial_clause[1][141] 	= partial_clause_prev[1][141] & 1'b1;
			partial_clause[1][142] 	= partial_clause_prev[1][142] & 1'b1;
			partial_clause[1][143] 	= partial_clause_prev[1][143] & 1'b1;
			partial_clause[1][144] 	= partial_clause_prev[1][144] & x[13];
			partial_clause[1][145] 	= partial_clause_prev[1][145] & 1'b1;
			partial_clause[1][146] 	= partial_clause_prev[1][146] & 1'b1;
			partial_clause[1][147] 	= partial_clause_prev[1][147] & 1'b1;
			partial_clause[1][148] 	= partial_clause_prev[1][148] & 1'b1;
			partial_clause[1][149] 	= partial_clause_prev[1][149] & 1'b1;
			partial_clause[1][150] 	= partial_clause_prev[1][150] & 1'b1;
			partial_clause[1][151] 	= partial_clause_prev[1][151] & 1'b1;
			partial_clause[1][152] 	= partial_clause_prev[1][152] & 1'b1;
			partial_clause[1][153] 	= partial_clause_prev[1][153] & x[43];
			partial_clause[1][154] 	= partial_clause_prev[1][154] & 1'b1;
			partial_clause[1][155] 	= partial_clause_prev[1][155] & 1'b1;
			partial_clause[1][156] 	= partial_clause_prev[1][156] & x[44];
			partial_clause[1][157] 	= partial_clause_prev[1][157] & 1'b1;
			partial_clause[1][158] 	= partial_clause_prev[1][158] & 1'b1;
			partial_clause[1][159] 	= partial_clause_prev[1][159] & 1'b1;
			partial_clause[1][160] 	= partial_clause_prev[1][160] & 1'b1;
			partial_clause[1][161] 	= partial_clause_prev[1][161] & 1'b1;
			partial_clause[1][162] 	= partial_clause_prev[1][162] & x[40];
			partial_clause[1][163] 	= partial_clause_prev[1][163] & 1'b1;
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & x[13];
			partial_clause[1][166] 	= partial_clause_prev[1][166] & 1'b1;
			partial_clause[1][167] 	= partial_clause_prev[1][167] & 1'b1;
			partial_clause[1][168] 	= partial_clause_prev[1][168] & 1'b1;
			partial_clause[1][169] 	= partial_clause_prev[1][169] & 1'b1;
			partial_clause[1][170] 	= partial_clause_prev[1][170] & 1'b1;
			partial_clause[1][171] 	= partial_clause_prev[1][171] & 1'b1;
			partial_clause[1][172] 	= partial_clause_prev[1][172] & 1'b1;
			partial_clause[1][173] 	= partial_clause_prev[1][173] & 1'b1;
			partial_clause[1][174] 	= partial_clause_prev[1][174] & 1'b1;
			partial_clause[1][175] 	= partial_clause_prev[1][175] & 1'b1;
			partial_clause[1][176] 	= partial_clause_prev[1][176] & 1'b1;
			partial_clause[1][177] 	= partial_clause_prev[1][177] & 1'b1;
			partial_clause[1][178] 	= partial_clause_prev[1][178] & 1'b1;
			partial_clause[1][179] 	= partial_clause_prev[1][179] & 1'b1;
			partial_clause[1][180] 	= partial_clause_prev[1][180] & 1'b1;
			partial_clause[1][181] 	= partial_clause_prev[1][181] & 1'b1;
			partial_clause[1][182] 	= partial_clause_prev[1][182] & 1'b1;
			partial_clause[1][183] 	= partial_clause_prev[1][183] & 1'b1;
			partial_clause[1][184] 	= partial_clause_prev[1][184] & 1'b1;
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & x[40];
			partial_clause[1][187] 	= partial_clause_prev[1][187] & 1'b1;
			partial_clause[1][188] 	= partial_clause_prev[1][188] & 1'b1;
			partial_clause[1][189] 	= partial_clause_prev[1][189] & 1'b1;
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & 1'b1;
			partial_clause[1][192] 	= partial_clause_prev[1][192] & 1'b1;
			partial_clause[1][193] 	= partial_clause_prev[1][193] & x[19];
			partial_clause[1][194] 	= partial_clause_prev[1][194] & 1'b1;
			partial_clause[1][195] 	= partial_clause_prev[1][195] & x[40];
			partial_clause[1][196] 	= partial_clause_prev[1][196] & 1'b1;
			partial_clause[1][197] 	= partial_clause_prev[1][197] & 1'b1;
			partial_clause[1][198] 	= partial_clause_prev[1][198] & 1'b1;
			partial_clause[1][199] 	= partial_clause_prev[1][199] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & x[3];
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & ~x[46];
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & ~x[44];
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & 1'b1;
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & x[17];
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			partial_clause[2][100] 	= partial_clause_prev[2][100] & 1'b1;
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & ~x[60];
			partial_clause[2][103] 	= partial_clause_prev[2][103] & 1'b1;
			partial_clause[2][104] 	= partial_clause_prev[2][104] & 1'b1;
			partial_clause[2][105] 	= partial_clause_prev[2][105] & 1'b1;
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & 1'b1;
			partial_clause[2][108] 	= partial_clause_prev[2][108] & 1'b1;
			partial_clause[2][109] 	= partial_clause_prev[2][109] & 1'b1;
			partial_clause[2][110] 	= partial_clause_prev[2][110] & 1'b1;
			partial_clause[2][111] 	= partial_clause_prev[2][111] & 1'b1;
			partial_clause[2][112] 	= partial_clause_prev[2][112] & 1'b1;
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & 1'b1;
			partial_clause[2][115] 	= partial_clause_prev[2][115] & 1'b1;
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & 1'b1;
			partial_clause[2][118] 	= partial_clause_prev[2][118] & 1'b1;
			partial_clause[2][119] 	= partial_clause_prev[2][119] & 1'b1;
			partial_clause[2][120] 	= partial_clause_prev[2][120] & 1'b1;
			partial_clause[2][121] 	= partial_clause_prev[2][121] & 1'b1;
			partial_clause[2][122] 	= partial_clause_prev[2][122] & 1'b1;
			partial_clause[2][123] 	= partial_clause_prev[2][123] & 1'b1;
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & 1'b1;
			partial_clause[2][126] 	= partial_clause_prev[2][126] & 1'b1;
			partial_clause[2][127] 	= partial_clause_prev[2][127] & 1'b1;
			partial_clause[2][128] 	= partial_clause_prev[2][128] & 1'b1;
			partial_clause[2][129] 	= partial_clause_prev[2][129] & 1'b1;
			partial_clause[2][130] 	= partial_clause_prev[2][130] & 1'b1;
			partial_clause[2][131] 	= partial_clause_prev[2][131] & 1'b1;
			partial_clause[2][132] 	= partial_clause_prev[2][132] & 1'b1;
			partial_clause[2][133] 	= partial_clause_prev[2][133] & 1'b1;
			partial_clause[2][134] 	= partial_clause_prev[2][134] & 1'b1;
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & 1'b1;
			partial_clause[2][137] 	= partial_clause_prev[2][137] & 1'b1;
			partial_clause[2][138] 	= partial_clause_prev[2][138] & 1'b1;
			partial_clause[2][139] 	= partial_clause_prev[2][139] & 1'b1;
			partial_clause[2][140] 	= partial_clause_prev[2][140] & 1'b1;
			partial_clause[2][141] 	= partial_clause_prev[2][141] & 1'b1;
			partial_clause[2][142] 	= partial_clause_prev[2][142] & 1'b1;
			partial_clause[2][143] 	= partial_clause_prev[2][143] & 1'b1;
			partial_clause[2][144] 	= partial_clause_prev[2][144] & 1'b1;
			partial_clause[2][145] 	= partial_clause_prev[2][145] & 1'b1;
			partial_clause[2][146] 	= partial_clause_prev[2][146] & 1'b1;
			partial_clause[2][147] 	= partial_clause_prev[2][147] & 1'b1;
			partial_clause[2][148] 	= partial_clause_prev[2][148] & 1'b1;
			partial_clause[2][149] 	= partial_clause_prev[2][149] & 1'b1;
			partial_clause[2][150] 	= partial_clause_prev[2][150] & 1'b1;
			partial_clause[2][151] 	= partial_clause_prev[2][151] & 1'b1;
			partial_clause[2][152] 	= partial_clause_prev[2][152] & 1'b1;
			partial_clause[2][153] 	= partial_clause_prev[2][153] & 1'b1;
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & 1'b1;
			partial_clause[2][156] 	= partial_clause_prev[2][156] & 1'b1;
			partial_clause[2][157] 	= partial_clause_prev[2][157] & 1'b1;
			partial_clause[2][158] 	= partial_clause_prev[2][158] & 1'b1;
			partial_clause[2][159] 	= partial_clause_prev[2][159] & 1'b1;
			partial_clause[2][160] 	= partial_clause_prev[2][160] & 1'b1;
			partial_clause[2][161] 	= partial_clause_prev[2][161] & 1'b1;
			partial_clause[2][162] 	= partial_clause_prev[2][162] & 1'b1;
			partial_clause[2][163] 	= partial_clause_prev[2][163] & 1'b1;
			partial_clause[2][164] 	= partial_clause_prev[2][164] & 1'b1;
			partial_clause[2][165] 	= partial_clause_prev[2][165] & 1'b1;
			partial_clause[2][166] 	= partial_clause_prev[2][166] & 1'b1;
			partial_clause[2][167] 	= partial_clause_prev[2][167] & 1'b1;
			partial_clause[2][168] 	= partial_clause_prev[2][168] & 1'b1;
			partial_clause[2][169] 	= partial_clause_prev[2][169] & 1'b1;
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & 1'b1;
			partial_clause[2][173] 	= partial_clause_prev[2][173] & 1'b1;
			partial_clause[2][174] 	= partial_clause_prev[2][174] & 1'b1;
			partial_clause[2][175] 	= partial_clause_prev[2][175] & x[63];
			partial_clause[2][176] 	= partial_clause_prev[2][176] & 1'b1;
			partial_clause[2][177] 	= partial_clause_prev[2][177] & 1'b1;
			partial_clause[2][178] 	= partial_clause_prev[2][178] & 1'b1;
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & 1'b1;
			partial_clause[2][181] 	= partial_clause_prev[2][181] & 1'b1;
			partial_clause[2][182] 	= partial_clause_prev[2][182] & 1'b1;
			partial_clause[2][183] 	= partial_clause_prev[2][183] & 1'b1;
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & 1'b1;
			partial_clause[2][186] 	= partial_clause_prev[2][186] & 1'b1;
			partial_clause[2][187] 	= partial_clause_prev[2][187] & 1'b1;
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & 1'b1;
			partial_clause[2][190] 	= partial_clause_prev[2][190] & 1'b1;
			partial_clause[2][191] 	= partial_clause_prev[2][191] & 1'b1;
			partial_clause[2][192] 	= partial_clause_prev[2][192] & 1'b1;
			partial_clause[2][193] 	= partial_clause_prev[2][193] & 1'b1;
			partial_clause[2][194] 	= partial_clause_prev[2][194] & 1'b1;
			partial_clause[2][195] 	= partial_clause_prev[2][195] & 1'b1;
			partial_clause[2][196] 	= partial_clause_prev[2][196] & 1'b1;
			partial_clause[2][197] 	= partial_clause_prev[2][197] & 1'b1;
			partial_clause[2][198] 	= partial_clause_prev[2][198] & 1'b1;
			partial_clause[2][199] 	= partial_clause_prev[2][199] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & ~x[43];
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & ~x[54];
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & x[8];
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & ~x[54];
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & ~x[27];
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & ~x[55];
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & x[16];
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & x[8];
			partial_clause[3][40] 	= partial_clause_prev[3][40] & ~x[39];
			partial_clause[3][41] 	= partial_clause_prev[3][41] & ~x[55];
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & ~x[45];
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[26];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & x[21];
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & x[48];
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & ~x[44];
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & x[10];
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			partial_clause[3][100] 	= partial_clause_prev[3][100] & 1'b1;
			partial_clause[3][101] 	= partial_clause_prev[3][101] & 1'b1;
			partial_clause[3][102] 	= partial_clause_prev[3][102] & 1'b1;
			partial_clause[3][103] 	= partial_clause_prev[3][103] & 1'b1;
			partial_clause[3][104] 	= partial_clause_prev[3][104] & 1'b1;
			partial_clause[3][105] 	= partial_clause_prev[3][105] & 1'b1;
			partial_clause[3][106] 	= partial_clause_prev[3][106] & 1'b1;
			partial_clause[3][107] 	= partial_clause_prev[3][107] & 1'b1;
			partial_clause[3][108] 	= partial_clause_prev[3][108] & 1'b1;
			partial_clause[3][109] 	= partial_clause_prev[3][109] & 1'b1;
			partial_clause[3][110] 	= partial_clause_prev[3][110] & 1'b1;
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & x[27];
			partial_clause[3][113] 	= partial_clause_prev[3][113] & 1'b1;
			partial_clause[3][114] 	= partial_clause_prev[3][114] & 1'b1;
			partial_clause[3][115] 	= partial_clause_prev[3][115] & ~x[12];
			partial_clause[3][116] 	= partial_clause_prev[3][116] & 1'b1;
			partial_clause[3][117] 	= partial_clause_prev[3][117] & 1'b1;
			partial_clause[3][118] 	= partial_clause_prev[3][118] & 1'b1;
			partial_clause[3][119] 	= partial_clause_prev[3][119] & 1'b1;
			partial_clause[3][120] 	= partial_clause_prev[3][120] & 1'b1;
			partial_clause[3][121] 	= partial_clause_prev[3][121] & 1'b1;
			partial_clause[3][122] 	= partial_clause_prev[3][122] & ~x[53];
			partial_clause[3][123] 	= partial_clause_prev[3][123] & 1'b1;
			partial_clause[3][124] 	= partial_clause_prev[3][124] & 1'b1;
			partial_clause[3][125] 	= partial_clause_prev[3][125] & 1'b1;
			partial_clause[3][126] 	= partial_clause_prev[3][126] & 1'b1;
			partial_clause[3][127] 	= partial_clause_prev[3][127] & 1'b1;
			partial_clause[3][128] 	= partial_clause_prev[3][128] & ~x[38];
			partial_clause[3][129] 	= partial_clause_prev[3][129] & 1'b1;
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & x[0];
			partial_clause[3][132] 	= partial_clause_prev[3][132] & 1'b1;
			partial_clause[3][133] 	= partial_clause_prev[3][133] & 1'b1;
			partial_clause[3][134] 	= partial_clause_prev[3][134] & 1'b1;
			partial_clause[3][135] 	= partial_clause_prev[3][135] & 1'b1;
			partial_clause[3][136] 	= partial_clause_prev[3][136] & 1'b1;
			partial_clause[3][137] 	= partial_clause_prev[3][137] & 1'b1;
			partial_clause[3][138] 	= partial_clause_prev[3][138] & 1'b1;
			partial_clause[3][139] 	= partial_clause_prev[3][139] & 1'b1;
			partial_clause[3][140] 	= partial_clause_prev[3][140] & 1'b1;
			partial_clause[3][141] 	= partial_clause_prev[3][141] & 1'b1;
			partial_clause[3][142] 	= partial_clause_prev[3][142] & 1'b1;
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & 1'b1;
			partial_clause[3][145] 	= partial_clause_prev[3][145] & ~x[14];
			partial_clause[3][146] 	= partial_clause_prev[3][146] & 1'b1;
			partial_clause[3][147] 	= partial_clause_prev[3][147] & 1'b1;
			partial_clause[3][148] 	= partial_clause_prev[3][148] & 1'b1;
			partial_clause[3][149] 	= partial_clause_prev[3][149] & ~x[19] & ~x[20];
			partial_clause[3][150] 	= partial_clause_prev[3][150] & 1'b1;
			partial_clause[3][151] 	= partial_clause_prev[3][151] & 1'b1;
			partial_clause[3][152] 	= partial_clause_prev[3][152] & 1'b1;
			partial_clause[3][153] 	= partial_clause_prev[3][153] & 1'b1;
			partial_clause[3][154] 	= partial_clause_prev[3][154] & 1'b1;
			partial_clause[3][155] 	= partial_clause_prev[3][155] & 1'b1;
			partial_clause[3][156] 	= partial_clause_prev[3][156] & 1'b1;
			partial_clause[3][157] 	= partial_clause_prev[3][157] & 1'b1;
			partial_clause[3][158] 	= partial_clause_prev[3][158] & 1'b1;
			partial_clause[3][159] 	= partial_clause_prev[3][159] & 1'b1;
			partial_clause[3][160] 	= partial_clause_prev[3][160] & 1'b1;
			partial_clause[3][161] 	= partial_clause_prev[3][161] & 1'b1;
			partial_clause[3][162] 	= partial_clause_prev[3][162] & 1'b1;
			partial_clause[3][163] 	= partial_clause_prev[3][163] & 1'b1;
			partial_clause[3][164] 	= partial_clause_prev[3][164] & 1'b1;
			partial_clause[3][165] 	= partial_clause_prev[3][165] & 1'b1;
			partial_clause[3][166] 	= partial_clause_prev[3][166] & 1'b1;
			partial_clause[3][167] 	= partial_clause_prev[3][167] & 1'b1;
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & 1'b1;
			partial_clause[3][170] 	= partial_clause_prev[3][170] & 1'b1;
			partial_clause[3][171] 	= partial_clause_prev[3][171] & 1'b1;
			partial_clause[3][172] 	= partial_clause_prev[3][172] & 1'b1;
			partial_clause[3][173] 	= partial_clause_prev[3][173] & ~x[16];
			partial_clause[3][174] 	= partial_clause_prev[3][174] & 1'b1;
			partial_clause[3][175] 	= partial_clause_prev[3][175] & 1'b1;
			partial_clause[3][176] 	= partial_clause_prev[3][176] & 1'b1;
			partial_clause[3][177] 	= partial_clause_prev[3][177] & 1'b1;
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & 1'b1;
			partial_clause[3][180] 	= partial_clause_prev[3][180] & ~x[7];
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & 1'b1;
			partial_clause[3][183] 	= partial_clause_prev[3][183] & 1'b1;
			partial_clause[3][184] 	= partial_clause_prev[3][184] & 1'b1;
			partial_clause[3][185] 	= partial_clause_prev[3][185] & 1'b1;
			partial_clause[3][186] 	= partial_clause_prev[3][186] & 1'b1;
			partial_clause[3][187] 	= partial_clause_prev[3][187] & 1'b1;
			partial_clause[3][188] 	= partial_clause_prev[3][188] & 1'b1;
			partial_clause[3][189] 	= partial_clause_prev[3][189] & 1'b1;
			partial_clause[3][190] 	= partial_clause_prev[3][190] & x[28];
			partial_clause[3][191] 	= partial_clause_prev[3][191] & 1'b1;
			partial_clause[3][192] 	= partial_clause_prev[3][192] & 1'b1;
			partial_clause[3][193] 	= partial_clause_prev[3][193] & 1'b1;
			partial_clause[3][194] 	= partial_clause_prev[3][194] & 1'b1;
			partial_clause[3][195] 	= partial_clause_prev[3][195] & 1'b1;
			partial_clause[3][196] 	= partial_clause_prev[3][196] & 1'b1;
			partial_clause[3][197] 	= partial_clause_prev[3][197] & 1'b1;
			partial_clause[3][198] 	= partial_clause_prev[3][198] & 1'b1;
			partial_clause[3][199] 	= partial_clause_prev[3][199] & ~x[15];
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & ~x[46];
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & ~x[47];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & ~x[44];
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & x[33];
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & ~x[18];
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & ~x[21] & ~x[48];
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & ~x[19];
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[47];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & ~x[13];
			partial_clause[4][35] 	= partial_clause_prev[4][35] & ~x[48];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & ~x[20];
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & ~x[19] & ~x[46];
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[45] & ~x[46];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & ~x[18];
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & ~x[44];
			partial_clause[4][53] 	= partial_clause_prev[4][53] & ~x[20];
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & ~x[46];
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & ~x[21];
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & ~x[17] & ~x[45];
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & ~x[19];
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & ~x[47];
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & ~x[20] & ~x[48];
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & x[58];
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			partial_clause[4][100] 	= partial_clause_prev[4][100] & 1'b1;
			partial_clause[4][101] 	= partial_clause_prev[4][101] & 1'b1;
			partial_clause[4][102] 	= partial_clause_prev[4][102] & x[19] & x[20] & x[44];
			partial_clause[4][103] 	= partial_clause_prev[4][103] & x[21];
			partial_clause[4][104] 	= partial_clause_prev[4][104] & 1'b1;
			partial_clause[4][105] 	= partial_clause_prev[4][105] & x[12];
			partial_clause[4][106] 	= partial_clause_prev[4][106] & x[20] & x[44];
			partial_clause[4][107] 	= partial_clause_prev[4][107] & 1'b1;
			partial_clause[4][108] 	= partial_clause_prev[4][108] & 1'b1;
			partial_clause[4][109] 	= partial_clause_prev[4][109] & x[47];
			partial_clause[4][110] 	= partial_clause_prev[4][110] & 1'b1;
			partial_clause[4][111] 	= partial_clause_prev[4][111] & 1'b1;
			partial_clause[4][112] 	= partial_clause_prev[4][112] & 1'b1;
			partial_clause[4][113] 	= partial_clause_prev[4][113] & 1'b1;
			partial_clause[4][114] 	= partial_clause_prev[4][114] & 1'b1;
			partial_clause[4][115] 	= partial_clause_prev[4][115] & 1'b1;
			partial_clause[4][116] 	= partial_clause_prev[4][116] & ~x[26];
			partial_clause[4][117] 	= partial_clause_prev[4][117] & 1'b1;
			partial_clause[4][118] 	= partial_clause_prev[4][118] & 1'b1;
			partial_clause[4][119] 	= partial_clause_prev[4][119] & 1'b1;
			partial_clause[4][120] 	= partial_clause_prev[4][120] & 1'b1;
			partial_clause[4][121] 	= partial_clause_prev[4][121] & 1'b1;
			partial_clause[4][122] 	= partial_clause_prev[4][122] & x[18];
			partial_clause[4][123] 	= partial_clause_prev[4][123] & 1'b1;
			partial_clause[4][124] 	= partial_clause_prev[4][124] & 1'b1;
			partial_clause[4][125] 	= partial_clause_prev[4][125] & 1'b1;
			partial_clause[4][126] 	= partial_clause_prev[4][126] & 1'b1;
			partial_clause[4][127] 	= partial_clause_prev[4][127] & 1'b1;
			partial_clause[4][128] 	= partial_clause_prev[4][128] & 1'b1;
			partial_clause[4][129] 	= partial_clause_prev[4][129] & 1'b1;
			partial_clause[4][130] 	= partial_clause_prev[4][130] & 1'b1;
			partial_clause[4][131] 	= partial_clause_prev[4][131] & x[18] & ~x[27];
			partial_clause[4][132] 	= partial_clause_prev[4][132] & 1'b1;
			partial_clause[4][133] 	= partial_clause_prev[4][133] & 1'b1;
			partial_clause[4][134] 	= partial_clause_prev[4][134] & 1'b1;
			partial_clause[4][135] 	= partial_clause_prev[4][135] & 1'b1;
			partial_clause[4][136] 	= partial_clause_prev[4][136] & 1'b1;
			partial_clause[4][137] 	= partial_clause_prev[4][137] & 1'b1;
			partial_clause[4][138] 	= partial_clause_prev[4][138] & 1'b1;
			partial_clause[4][139] 	= partial_clause_prev[4][139] & 1'b1;
			partial_clause[4][140] 	= partial_clause_prev[4][140] & 1'b1;
			partial_clause[4][141] 	= partial_clause_prev[4][141] & 1'b1;
			partial_clause[4][142] 	= partial_clause_prev[4][142] & 1'b1;
			partial_clause[4][143] 	= partial_clause_prev[4][143] & 1'b1;
			partial_clause[4][144] 	= partial_clause_prev[4][144] & x[17] & x[18] & x[20];
			partial_clause[4][145] 	= partial_clause_prev[4][145] & 1'b1;
			partial_clause[4][146] 	= partial_clause_prev[4][146] & 1'b1;
			partial_clause[4][147] 	= partial_clause_prev[4][147] & 1'b1;
			partial_clause[4][148] 	= partial_clause_prev[4][148] & x[13];
			partial_clause[4][149] 	= partial_clause_prev[4][149] & 1'b1;
			partial_clause[4][150] 	= partial_clause_prev[4][150] & 1'b1;
			partial_clause[4][151] 	= partial_clause_prev[4][151] & x[16];
			partial_clause[4][152] 	= partial_clause_prev[4][152] & 1'b1;
			partial_clause[4][153] 	= partial_clause_prev[4][153] & 1'b1;
			partial_clause[4][154] 	= partial_clause_prev[4][154] & 1'b1;
			partial_clause[4][155] 	= partial_clause_prev[4][155] & x[20] & x[21];
			partial_clause[4][156] 	= partial_clause_prev[4][156] & 1'b1;
			partial_clause[4][157] 	= partial_clause_prev[4][157] & x[45] & x[48];
			partial_clause[4][158] 	= partial_clause_prev[4][158] & 1'b1;
			partial_clause[4][159] 	= partial_clause_prev[4][159] & 1'b1;
			partial_clause[4][160] 	= partial_clause_prev[4][160] & x[18] & x[19] & x[20];
			partial_clause[4][161] 	= partial_clause_prev[4][161] & 1'b1;
			partial_clause[4][162] 	= partial_clause_prev[4][162] & x[22] & x[46];
			partial_clause[4][163] 	= partial_clause_prev[4][163] & 1'b1;
			partial_clause[4][164] 	= partial_clause_prev[4][164] & x[46] & x[48];
			partial_clause[4][165] 	= partial_clause_prev[4][165] & x[43];
			partial_clause[4][166] 	= partial_clause_prev[4][166] & 1'b1;
			partial_clause[4][167] 	= partial_clause_prev[4][167] & 1'b1;
			partial_clause[4][168] 	= partial_clause_prev[4][168] & 1'b1;
			partial_clause[4][169] 	= partial_clause_prev[4][169] & 1'b1;
			partial_clause[4][170] 	= partial_clause_prev[4][170] & 1'b1;
			partial_clause[4][171] 	= partial_clause_prev[4][171] & 1'b1;
			partial_clause[4][172] 	= partial_clause_prev[4][172] & 1'b1;
			partial_clause[4][173] 	= partial_clause_prev[4][173] & 1'b1;
			partial_clause[4][174] 	= partial_clause_prev[4][174] & x[16] & x[17];
			partial_clause[4][175] 	= partial_clause_prev[4][175] & 1'b1;
			partial_clause[4][176] 	= partial_clause_prev[4][176] & 1'b1;
			partial_clause[4][177] 	= partial_clause_prev[4][177] & 1'b1;
			partial_clause[4][178] 	= partial_clause_prev[4][178] & 1'b1;
			partial_clause[4][179] 	= partial_clause_prev[4][179] & 1'b1;
			partial_clause[4][180] 	= partial_clause_prev[4][180] & 1'b1;
			partial_clause[4][181] 	= partial_clause_prev[4][181] & 1'b1;
			partial_clause[4][182] 	= partial_clause_prev[4][182] & x[21] & x[23];
			partial_clause[4][183] 	= partial_clause_prev[4][183] & 1'b1;
			partial_clause[4][184] 	= partial_clause_prev[4][184] & 1'b1;
			partial_clause[4][185] 	= partial_clause_prev[4][185] & 1'b1;
			partial_clause[4][186] 	= partial_clause_prev[4][186] & 1'b1;
			partial_clause[4][187] 	= partial_clause_prev[4][187] & x[16];
			partial_clause[4][188] 	= partial_clause_prev[4][188] & 1'b1;
			partial_clause[4][189] 	= partial_clause_prev[4][189] & 1'b1;
			partial_clause[4][190] 	= partial_clause_prev[4][190] & 1'b1;
			partial_clause[4][191] 	= partial_clause_prev[4][191] & 1'b1;
			partial_clause[4][192] 	= partial_clause_prev[4][192] & 1'b1;
			partial_clause[4][193] 	= partial_clause_prev[4][193] & 1'b1;
			partial_clause[4][194] 	= partial_clause_prev[4][194] & 1'b1;
			partial_clause[4][195] 	= partial_clause_prev[4][195] & x[46] & x[47];
			partial_clause[4][196] 	= partial_clause_prev[4][196] & 1'b1;
			partial_clause[4][197] 	= partial_clause_prev[4][197] & x[41];
			partial_clause[4][198] 	= partial_clause_prev[4][198] & ~x[27];
			partial_clause[4][199] 	= partial_clause_prev[4][199] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & x[43];
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & x[28];
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & ~x[48];
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & x[50];
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & ~x[10];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & ~x[47] & ~x[49] & ~x[51] & ~x[53];
			partial_clause[5][29] 	= partial_clause_prev[5][29] & x[25];
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & x[0];
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & ~x[53];
			partial_clause[5][41] 	= partial_clause_prev[5][41] & x[57];
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & x[57];
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & x[40];
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & x[52];
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & x[22];
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & ~x[21];
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & x[21] & x[23];
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & x[24];
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & ~x[19] & ~x[20] & ~x[21] & ~x[23];
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & x[0];
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & ~x[53];
			partial_clause[5][82] 	= partial_clause_prev[5][82] & x[52];
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & x[27];
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & x[21];
			partial_clause[5][96] 	= partial_clause_prev[5][96] & x[29];
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			partial_clause[5][100] 	= partial_clause_prev[5][100] & x[8];
			partial_clause[5][101] 	= partial_clause_prev[5][101] & 1'b1;
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & 1'b1;
			partial_clause[5][104] 	= partial_clause_prev[5][104] & 1'b1;
			partial_clause[5][105] 	= partial_clause_prev[5][105] & 1'b1;
			partial_clause[5][106] 	= partial_clause_prev[5][106] & 1'b1;
			partial_clause[5][107] 	= partial_clause_prev[5][107] & 1'b1;
			partial_clause[5][108] 	= partial_clause_prev[5][108] & 1'b1;
			partial_clause[5][109] 	= partial_clause_prev[5][109] & ~x[54];
			partial_clause[5][110] 	= partial_clause_prev[5][110] & ~x[54];
			partial_clause[5][111] 	= partial_clause_prev[5][111] & 1'b1;
			partial_clause[5][112] 	= partial_clause_prev[5][112] & 1'b1;
			partial_clause[5][113] 	= partial_clause_prev[5][113] & 1'b1;
			partial_clause[5][114] 	= partial_clause_prev[5][114] & 1'b1;
			partial_clause[5][115] 	= partial_clause_prev[5][115] & 1'b1;
			partial_clause[5][116] 	= partial_clause_prev[5][116] & 1'b1;
			partial_clause[5][117] 	= partial_clause_prev[5][117] & x[24];
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & 1'b1;
			partial_clause[5][120] 	= partial_clause_prev[5][120] & 1'b1;
			partial_clause[5][121] 	= partial_clause_prev[5][121] & 1'b1;
			partial_clause[5][122] 	= partial_clause_prev[5][122] & 1'b1;
			partial_clause[5][123] 	= partial_clause_prev[5][123] & 1'b1;
			partial_clause[5][124] 	= partial_clause_prev[5][124] & 1'b1;
			partial_clause[5][125] 	= partial_clause_prev[5][125] & 1'b1;
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & 1'b1;
			partial_clause[5][128] 	= partial_clause_prev[5][128] & 1'b1;
			partial_clause[5][129] 	= partial_clause_prev[5][129] & 1'b1;
			partial_clause[5][130] 	= partial_clause_prev[5][130] & 1'b1;
			partial_clause[5][131] 	= partial_clause_prev[5][131] & 1'b1;
			partial_clause[5][132] 	= partial_clause_prev[5][132] & ~x[26];
			partial_clause[5][133] 	= partial_clause_prev[5][133] & 1'b1;
			partial_clause[5][134] 	= partial_clause_prev[5][134] & 1'b1;
			partial_clause[5][135] 	= partial_clause_prev[5][135] & 1'b1;
			partial_clause[5][136] 	= partial_clause_prev[5][136] & 1'b1;
			partial_clause[5][137] 	= partial_clause_prev[5][137] & 1'b1;
			partial_clause[5][138] 	= partial_clause_prev[5][138] & 1'b1;
			partial_clause[5][139] 	= partial_clause_prev[5][139] & 1'b1;
			partial_clause[5][140] 	= partial_clause_prev[5][140] & 1'b1;
			partial_clause[5][141] 	= partial_clause_prev[5][141] & 1'b1;
			partial_clause[5][142] 	= partial_clause_prev[5][142] & 1'b1;
			partial_clause[5][143] 	= partial_clause_prev[5][143] & 1'b1;
			partial_clause[5][144] 	= partial_clause_prev[5][144] & 1'b1;
			partial_clause[5][145] 	= partial_clause_prev[5][145] & 1'b1;
			partial_clause[5][146] 	= partial_clause_prev[5][146] & 1'b1;
			partial_clause[5][147] 	= partial_clause_prev[5][147] & 1'b1;
			partial_clause[5][148] 	= partial_clause_prev[5][148] & 1'b1;
			partial_clause[5][149] 	= partial_clause_prev[5][149] & 1'b1;
			partial_clause[5][150] 	= partial_clause_prev[5][150] & 1'b1;
			partial_clause[5][151] 	= partial_clause_prev[5][151] & 1'b1;
			partial_clause[5][152] 	= partial_clause_prev[5][152] & ~x[26];
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & 1'b1;
			partial_clause[5][155] 	= partial_clause_prev[5][155] & 1'b1;
			partial_clause[5][156] 	= partial_clause_prev[5][156] & 1'b1;
			partial_clause[5][157] 	= partial_clause_prev[5][157] & ~x[0];
			partial_clause[5][158] 	= partial_clause_prev[5][158] & 1'b1;
			partial_clause[5][159] 	= partial_clause_prev[5][159] & 1'b1;
			partial_clause[5][160] 	= partial_clause_prev[5][160] & 1'b1;
			partial_clause[5][161] 	= partial_clause_prev[5][161] & ~x[57];
			partial_clause[5][162] 	= partial_clause_prev[5][162] & 1'b1;
			partial_clause[5][163] 	= partial_clause_prev[5][163] & 1'b1;
			partial_clause[5][164] 	= partial_clause_prev[5][164] & ~x[0] & ~x[27] & ~x[28] & ~x[55];
			partial_clause[5][165] 	= partial_clause_prev[5][165] & 1'b1;
			partial_clause[5][166] 	= partial_clause_prev[5][166] & 1'b1;
			partial_clause[5][167] 	= partial_clause_prev[5][167] & 1'b1;
			partial_clause[5][168] 	= partial_clause_prev[5][168] & 1'b1;
			partial_clause[5][169] 	= partial_clause_prev[5][169] & 1'b1;
			partial_clause[5][170] 	= partial_clause_prev[5][170] & 1'b1;
			partial_clause[5][171] 	= partial_clause_prev[5][171] & 1'b1;
			partial_clause[5][172] 	= partial_clause_prev[5][172] & 1'b1;
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & 1'b1;
			partial_clause[5][175] 	= partial_clause_prev[5][175] & 1'b1;
			partial_clause[5][176] 	= partial_clause_prev[5][176] & 1'b1;
			partial_clause[5][177] 	= partial_clause_prev[5][177] & 1'b1;
			partial_clause[5][178] 	= partial_clause_prev[5][178] & x[8];
			partial_clause[5][179] 	= partial_clause_prev[5][179] & ~x[55];
			partial_clause[5][180] 	= partial_clause_prev[5][180] & ~x[54];
			partial_clause[5][181] 	= partial_clause_prev[5][181] & ~x[26];
			partial_clause[5][182] 	= partial_clause_prev[5][182] & 1'b1;
			partial_clause[5][183] 	= partial_clause_prev[5][183] & 1'b1;
			partial_clause[5][184] 	= partial_clause_prev[5][184] & 1'b1;
			partial_clause[5][185] 	= partial_clause_prev[5][185] & 1'b1;
			partial_clause[5][186] 	= partial_clause_prev[5][186] & ~x[26] & ~x[55];
			partial_clause[5][187] 	= partial_clause_prev[5][187] & ~x[28];
			partial_clause[5][188] 	= partial_clause_prev[5][188] & 1'b1;
			partial_clause[5][189] 	= partial_clause_prev[5][189] & 1'b1;
			partial_clause[5][190] 	= partial_clause_prev[5][190] & 1'b1;
			partial_clause[5][191] 	= partial_clause_prev[5][191] & 1'b1;
			partial_clause[5][192] 	= partial_clause_prev[5][192] & 1'b1;
			partial_clause[5][193] 	= partial_clause_prev[5][193] & 1'b1;
			partial_clause[5][194] 	= partial_clause_prev[5][194] & 1'b1;
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & 1'b1;
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & 1'b1;
			partial_clause[5][199] 	= partial_clause_prev[5][199] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & ~x[44] & ~x[55];
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & ~x[23] & ~x[24] & ~x[48];
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & ~x[45];
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & ~x[18];
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & ~x[20] & ~x[22] & ~x[23] & ~x[55];
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & ~x[16];
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & ~x[22] & ~x[25] & ~x[26] & ~x[48];
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & ~x[12] & ~x[23];
			partial_clause[6][46] 	= partial_clause_prev[6][46] & ~x[13];
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & ~x[25] & ~x[50];
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & x[31];
			partial_clause[6][52] 	= partial_clause_prev[6][52] & ~x[21] & ~x[53];
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & ~x[25] & ~x[48] & ~x[50];
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & ~x[12];
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & ~x[21] & ~x[25];
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & ~x[19];
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & ~x[45];
			partial_clause[6][76] 	= partial_clause_prev[6][76] & ~x[43] & ~x[53];
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & ~x[22] & ~x[47];
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & ~x[44];
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & ~x[19];
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & ~x[22];
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & ~x[50];
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & ~x[19];
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & ~x[19] & ~x[26] & ~x[46];
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			partial_clause[6][100] 	= partial_clause_prev[6][100] & 1'b1;
			partial_clause[6][101] 	= partial_clause_prev[6][101] & 1'b1;
			partial_clause[6][102] 	= partial_clause_prev[6][102] & x[50];
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & 1'b1;
			partial_clause[6][105] 	= partial_clause_prev[6][105] & 1'b1;
			partial_clause[6][106] 	= partial_clause_prev[6][106] & 1'b1;
			partial_clause[6][107] 	= partial_clause_prev[6][107] & ~x[52];
			partial_clause[6][108] 	= partial_clause_prev[6][108] & 1'b1;
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & x[50];
			partial_clause[6][111] 	= partial_clause_prev[6][111] & 1'b1;
			partial_clause[6][112] 	= partial_clause_prev[6][112] & 1'b1;
			partial_clause[6][113] 	= partial_clause_prev[6][113] & 1'b1;
			partial_clause[6][114] 	= partial_clause_prev[6][114] & 1'b1;
			partial_clause[6][115] 	= partial_clause_prev[6][115] & x[46];
			partial_clause[6][116] 	= partial_clause_prev[6][116] & 1'b1;
			partial_clause[6][117] 	= partial_clause_prev[6][117] & 1'b1;
			partial_clause[6][118] 	= partial_clause_prev[6][118] & ~x[35];
			partial_clause[6][119] 	= partial_clause_prev[6][119] & 1'b1;
			partial_clause[6][120] 	= partial_clause_prev[6][120] & x[47];
			partial_clause[6][121] 	= partial_clause_prev[6][121] & 1'b1;
			partial_clause[6][122] 	= partial_clause_prev[6][122] & 1'b1;
			partial_clause[6][123] 	= partial_clause_prev[6][123] & 1'b1;
			partial_clause[6][124] 	= partial_clause_prev[6][124] & 1'b1;
			partial_clause[6][125] 	= partial_clause_prev[6][125] & 1'b1;
			partial_clause[6][126] 	= partial_clause_prev[6][126] & 1'b1;
			partial_clause[6][127] 	= partial_clause_prev[6][127] & 1'b1;
			partial_clause[6][128] 	= partial_clause_prev[6][128] & 1'b1;
			partial_clause[6][129] 	= partial_clause_prev[6][129] & 1'b1;
			partial_clause[6][130] 	= partial_clause_prev[6][130] & 1'b1;
			partial_clause[6][131] 	= partial_clause_prev[6][131] & x[52];
			partial_clause[6][132] 	= partial_clause_prev[6][132] & 1'b1;
			partial_clause[6][133] 	= partial_clause_prev[6][133] & x[14];
			partial_clause[6][134] 	= partial_clause_prev[6][134] & 1'b1;
			partial_clause[6][135] 	= partial_clause_prev[6][135] & 1'b1;
			partial_clause[6][136] 	= partial_clause_prev[6][136] & x[22];
			partial_clause[6][137] 	= partial_clause_prev[6][137] & 1'b1;
			partial_clause[6][138] 	= partial_clause_prev[6][138] & 1'b1;
			partial_clause[6][139] 	= partial_clause_prev[6][139] & x[48];
			partial_clause[6][140] 	= partial_clause_prev[6][140] & 1'b1;
			partial_clause[6][141] 	= partial_clause_prev[6][141] & 1'b1;
			partial_clause[6][142] 	= partial_clause_prev[6][142] & 1'b1;
			partial_clause[6][143] 	= partial_clause_prev[6][143] & x[48];
			partial_clause[6][144] 	= partial_clause_prev[6][144] & 1'b1;
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & x[51];
			partial_clause[6][147] 	= partial_clause_prev[6][147] & 1'b1;
			partial_clause[6][148] 	= partial_clause_prev[6][148] & 1'b1;
			partial_clause[6][149] 	= partial_clause_prev[6][149] & 1'b1;
			partial_clause[6][150] 	= partial_clause_prev[6][150] & 1'b1;
			partial_clause[6][151] 	= partial_clause_prev[6][151] & x[50];
			partial_clause[6][152] 	= partial_clause_prev[6][152] & 1'b1;
			partial_clause[6][153] 	= partial_clause_prev[6][153] & x[21];
			partial_clause[6][154] 	= partial_clause_prev[6][154] & 1'b1;
			partial_clause[6][155] 	= partial_clause_prev[6][155] & 1'b1;
			partial_clause[6][156] 	= partial_clause_prev[6][156] & x[49];
			partial_clause[6][157] 	= partial_clause_prev[6][157] & 1'b1;
			partial_clause[6][158] 	= partial_clause_prev[6][158] & 1'b1;
			partial_clause[6][159] 	= partial_clause_prev[6][159] & 1'b1;
			partial_clause[6][160] 	= partial_clause_prev[6][160] & 1'b1;
			partial_clause[6][161] 	= partial_clause_prev[6][161] & 1'b1;
			partial_clause[6][162] 	= partial_clause_prev[6][162] & 1'b1;
			partial_clause[6][163] 	= partial_clause_prev[6][163] & 1'b1;
			partial_clause[6][164] 	= partial_clause_prev[6][164] & 1'b1;
			partial_clause[6][165] 	= partial_clause_prev[6][165] & 1'b1;
			partial_clause[6][166] 	= partial_clause_prev[6][166] & x[52];
			partial_clause[6][167] 	= partial_clause_prev[6][167] & x[17];
			partial_clause[6][168] 	= partial_clause_prev[6][168] & x[19];
			partial_clause[6][169] 	= partial_clause_prev[6][169] & 1'b1;
			partial_clause[6][170] 	= partial_clause_prev[6][170] & 1'b1;
			partial_clause[6][171] 	= partial_clause_prev[6][171] & 1'b1;
			partial_clause[6][172] 	= partial_clause_prev[6][172] & 1'b1;
			partial_clause[6][173] 	= partial_clause_prev[6][173] & 1'b1;
			partial_clause[6][174] 	= partial_clause_prev[6][174] & 1'b1;
			partial_clause[6][175] 	= partial_clause_prev[6][175] & x[26];
			partial_clause[6][176] 	= partial_clause_prev[6][176] & 1'b1;
			partial_clause[6][177] 	= partial_clause_prev[6][177] & 1'b1;
			partial_clause[6][178] 	= partial_clause_prev[6][178] & 1'b1;
			partial_clause[6][179] 	= partial_clause_prev[6][179] & 1'b1;
			partial_clause[6][180] 	= partial_clause_prev[6][180] & 1'b1;
			partial_clause[6][181] 	= partial_clause_prev[6][181] & 1'b1;
			partial_clause[6][182] 	= partial_clause_prev[6][182] & 1'b1;
			partial_clause[6][183] 	= partial_clause_prev[6][183] & 1'b1;
			partial_clause[6][184] 	= partial_clause_prev[6][184] & x[54];
			partial_clause[6][185] 	= partial_clause_prev[6][185] & 1'b1;
			partial_clause[6][186] 	= partial_clause_prev[6][186] & 1'b1;
			partial_clause[6][187] 	= partial_clause_prev[6][187] & 1'b1;
			partial_clause[6][188] 	= partial_clause_prev[6][188] & 1'b1;
			partial_clause[6][189] 	= partial_clause_prev[6][189] & 1'b1;
			partial_clause[6][190] 	= partial_clause_prev[6][190] & 1'b1;
			partial_clause[6][191] 	= partial_clause_prev[6][191] & x[54];
			partial_clause[6][192] 	= partial_clause_prev[6][192] & 1'b1;
			partial_clause[6][193] 	= partial_clause_prev[6][193] & 1'b1;
			partial_clause[6][194] 	= partial_clause_prev[6][194] & 1'b1;
			partial_clause[6][195] 	= partial_clause_prev[6][195] & 1'b1;
			partial_clause[6][196] 	= partial_clause_prev[6][196] & 1'b1;
			partial_clause[6][197] 	= partial_clause_prev[6][197] & 1'b1;
			partial_clause[6][198] 	= partial_clause_prev[6][198] & x[26];
			partial_clause[6][199] 	= partial_clause_prev[6][199] & x[25];
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & x[50];
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & x[46] & x[49];
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & x[36];
			partial_clause[7][26] 	= partial_clause_prev[7][26] & x[31];
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & ~x[20];
			partial_clause[7][31] 	= partial_clause_prev[7][31] & x[45];
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & x[3];
			partial_clause[7][37] 	= partial_clause_prev[7][37] & ~x[18];
			partial_clause[7][38] 	= partial_clause_prev[7][38] & x[43];
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & x[43] & x[46];
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & x[16] & x[19] & x[49];
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & x[41];
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & x[40] & x[44];
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & x[12];
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & x[14];
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			partial_clause[7][100] 	= partial_clause_prev[7][100] & ~x[14];
			partial_clause[7][101] 	= partial_clause_prev[7][101] & 1'b1;
			partial_clause[7][102] 	= partial_clause_prev[7][102] & 1'b1;
			partial_clause[7][103] 	= partial_clause_prev[7][103] & 1'b1;
			partial_clause[7][104] 	= partial_clause_prev[7][104] & 1'b1;
			partial_clause[7][105] 	= partial_clause_prev[7][105] & ~x[46];
			partial_clause[7][106] 	= partial_clause_prev[7][106] & 1'b1;
			partial_clause[7][107] 	= partial_clause_prev[7][107] & 1'b1;
			partial_clause[7][108] 	= partial_clause_prev[7][108] & ~x[44];
			partial_clause[7][109] 	= partial_clause_prev[7][109] & ~x[14] & ~x[15] & ~x[43];
			partial_clause[7][110] 	= partial_clause_prev[7][110] & 1'b1;
			partial_clause[7][111] 	= partial_clause_prev[7][111] & 1'b1;
			partial_clause[7][112] 	= partial_clause_prev[7][112] & 1'b1;
			partial_clause[7][113] 	= partial_clause_prev[7][113] & 1'b1;
			partial_clause[7][114] 	= partial_clause_prev[7][114] & 1'b1;
			partial_clause[7][115] 	= partial_clause_prev[7][115] & 1'b1;
			partial_clause[7][116] 	= partial_clause_prev[7][116] & 1'b1;
			partial_clause[7][117] 	= partial_clause_prev[7][117] & 1'b1;
			partial_clause[7][118] 	= partial_clause_prev[7][118] & x[0];
			partial_clause[7][119] 	= partial_clause_prev[7][119] & 1'b1;
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & 1'b1;
			partial_clause[7][123] 	= partial_clause_prev[7][123] & 1'b1;
			partial_clause[7][124] 	= partial_clause_prev[7][124] & 1'b1;
			partial_clause[7][125] 	= partial_clause_prev[7][125] & 1'b1;
			partial_clause[7][126] 	= partial_clause_prev[7][126] & 1'b1;
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & 1'b1;
			partial_clause[7][129] 	= partial_clause_prev[7][129] & ~x[11] & ~x[39];
			partial_clause[7][130] 	= partial_clause_prev[7][130] & ~x[48] & ~x[49];
			partial_clause[7][131] 	= partial_clause_prev[7][131] & 1'b1;
			partial_clause[7][132] 	= partial_clause_prev[7][132] & 1'b1;
			partial_clause[7][133] 	= partial_clause_prev[7][133] & 1'b1;
			partial_clause[7][134] 	= partial_clause_prev[7][134] & 1'b1;
			partial_clause[7][135] 	= partial_clause_prev[7][135] & 1'b1;
			partial_clause[7][136] 	= partial_clause_prev[7][136] & 1'b1;
			partial_clause[7][137] 	= partial_clause_prev[7][137] & ~x[14] & ~x[41];
			partial_clause[7][138] 	= partial_clause_prev[7][138] & 1'b1;
			partial_clause[7][139] 	= partial_clause_prev[7][139] & 1'b1;
			partial_clause[7][140] 	= partial_clause_prev[7][140] & ~x[39];
			partial_clause[7][141] 	= partial_clause_prev[7][141] & ~x[15] & ~x[41] & ~x[42];
			partial_clause[7][142] 	= partial_clause_prev[7][142] & 1'b1;
			partial_clause[7][143] 	= partial_clause_prev[7][143] & 1'b1;
			partial_clause[7][144] 	= partial_clause_prev[7][144] & 1'b1;
			partial_clause[7][145] 	= partial_clause_prev[7][145] & 1'b1;
			partial_clause[7][146] 	= partial_clause_prev[7][146] & 1'b1;
			partial_clause[7][147] 	= partial_clause_prev[7][147] & 1'b1;
			partial_clause[7][148] 	= partial_clause_prev[7][148] & 1'b1;
			partial_clause[7][149] 	= partial_clause_prev[7][149] & 1'b1;
			partial_clause[7][150] 	= partial_clause_prev[7][150] & 1'b1;
			partial_clause[7][151] 	= partial_clause_prev[7][151] & 1'b1;
			partial_clause[7][152] 	= partial_clause_prev[7][152] & 1'b1;
			partial_clause[7][153] 	= partial_clause_prev[7][153] & 1'b1;
			partial_clause[7][154] 	= partial_clause_prev[7][154] & 1'b1;
			partial_clause[7][155] 	= partial_clause_prev[7][155] & 1'b1;
			partial_clause[7][156] 	= partial_clause_prev[7][156] & 1'b1;
			partial_clause[7][157] 	= partial_clause_prev[7][157] & 1'b1;
			partial_clause[7][158] 	= partial_clause_prev[7][158] & 1'b1;
			partial_clause[7][159] 	= partial_clause_prev[7][159] & 1'b1;
			partial_clause[7][160] 	= partial_clause_prev[7][160] & 1'b1;
			partial_clause[7][161] 	= partial_clause_prev[7][161] & 1'b1;
			partial_clause[7][162] 	= partial_clause_prev[7][162] & 1'b1;
			partial_clause[7][163] 	= partial_clause_prev[7][163] & 1'b1;
			partial_clause[7][164] 	= partial_clause_prev[7][164] & 1'b1;
			partial_clause[7][165] 	= partial_clause_prev[7][165] & 1'b1;
			partial_clause[7][166] 	= partial_clause_prev[7][166] & 1'b1;
			partial_clause[7][167] 	= partial_clause_prev[7][167] & 1'b1;
			partial_clause[7][168] 	= partial_clause_prev[7][168] & 1'b1;
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & 1'b1;
			partial_clause[7][171] 	= partial_clause_prev[7][171] & 1'b1;
			partial_clause[7][172] 	= partial_clause_prev[7][172] & 1'b1;
			partial_clause[7][173] 	= partial_clause_prev[7][173] & 1'b1;
			partial_clause[7][174] 	= partial_clause_prev[7][174] & 1'b1;
			partial_clause[7][175] 	= partial_clause_prev[7][175] & 1'b1;
			partial_clause[7][176] 	= partial_clause_prev[7][176] & 1'b1;
			partial_clause[7][177] 	= partial_clause_prev[7][177] & 1'b1;
			partial_clause[7][178] 	= partial_clause_prev[7][178] & 1'b1;
			partial_clause[7][179] 	= partial_clause_prev[7][179] & 1'b1;
			partial_clause[7][180] 	= partial_clause_prev[7][180] & 1'b1;
			partial_clause[7][181] 	= partial_clause_prev[7][181] & 1'b1;
			partial_clause[7][182] 	= partial_clause_prev[7][182] & 1'b1;
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & 1'b1;
			partial_clause[7][185] 	= partial_clause_prev[7][185] & 1'b1;
			partial_clause[7][186] 	= partial_clause_prev[7][186] & 1'b1;
			partial_clause[7][187] 	= partial_clause_prev[7][187] & 1'b1;
			partial_clause[7][188] 	= partial_clause_prev[7][188] & 1'b1;
			partial_clause[7][189] 	= partial_clause_prev[7][189] & 1'b1;
			partial_clause[7][190] 	= partial_clause_prev[7][190] & 1'b1;
			partial_clause[7][191] 	= partial_clause_prev[7][191] & 1'b1;
			partial_clause[7][192] 	= partial_clause_prev[7][192] & 1'b1;
			partial_clause[7][193] 	= partial_clause_prev[7][193] & ~x[41];
			partial_clause[7][194] 	= partial_clause_prev[7][194] & 1'b1;
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & 1'b1;
			partial_clause[7][197] 	= partial_clause_prev[7][197] & 1'b1;
			partial_clause[7][198] 	= partial_clause_prev[7][198] & ~x[16] & ~x[43];
			partial_clause[7][199] 	= partial_clause_prev[7][199] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & ~x[11];
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & ~x[19];
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & x[19];
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & ~x[46];
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & ~x[10];
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & ~x[11];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			partial_clause[8][100] 	= partial_clause_prev[8][100] & 1'b1;
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & ~x[15];
			partial_clause[8][103] 	= partial_clause_prev[8][103] & 1'b1;
			partial_clause[8][104] 	= partial_clause_prev[8][104] & 1'b1;
			partial_clause[8][105] 	= partial_clause_prev[8][105] & 1'b1;
			partial_clause[8][106] 	= partial_clause_prev[8][106] & 1'b1;
			partial_clause[8][107] 	= partial_clause_prev[8][107] & 1'b1;
			partial_clause[8][108] 	= partial_clause_prev[8][108] & 1'b1;
			partial_clause[8][109] 	= partial_clause_prev[8][109] & 1'b1;
			partial_clause[8][110] 	= partial_clause_prev[8][110] & 1'b1;
			partial_clause[8][111] 	= partial_clause_prev[8][111] & 1'b1;
			partial_clause[8][112] 	= partial_clause_prev[8][112] & 1'b1;
			partial_clause[8][113] 	= partial_clause_prev[8][113] & 1'b1;
			partial_clause[8][114] 	= partial_clause_prev[8][114] & 1'b1;
			partial_clause[8][115] 	= partial_clause_prev[8][115] & 1'b1;
			partial_clause[8][116] 	= partial_clause_prev[8][116] & 1'b1;
			partial_clause[8][117] 	= partial_clause_prev[8][117] & 1'b1;
			partial_clause[8][118] 	= partial_clause_prev[8][118] & 1'b1;
			partial_clause[8][119] 	= partial_clause_prev[8][119] & 1'b1;
			partial_clause[8][120] 	= partial_clause_prev[8][120] & 1'b1;
			partial_clause[8][121] 	= partial_clause_prev[8][121] & 1'b1;
			partial_clause[8][122] 	= partial_clause_prev[8][122] & x[62];
			partial_clause[8][123] 	= partial_clause_prev[8][123] & 1'b1;
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & 1'b1;
			partial_clause[8][126] 	= partial_clause_prev[8][126] & 1'b1;
			partial_clause[8][127] 	= partial_clause_prev[8][127] & 1'b1;
			partial_clause[8][128] 	= partial_clause_prev[8][128] & 1'b1;
			partial_clause[8][129] 	= partial_clause_prev[8][129] & 1'b1;
			partial_clause[8][130] 	= partial_clause_prev[8][130] & 1'b1;
			partial_clause[8][131] 	= partial_clause_prev[8][131] & 1'b1;
			partial_clause[8][132] 	= partial_clause_prev[8][132] & 1'b1;
			partial_clause[8][133] 	= partial_clause_prev[8][133] & 1'b1;
			partial_clause[8][134] 	= partial_clause_prev[8][134] & 1'b1;
			partial_clause[8][135] 	= partial_clause_prev[8][135] & ~x[55];
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & 1'b1;
			partial_clause[8][138] 	= partial_clause_prev[8][138] & 1'b1;
			partial_clause[8][139] 	= partial_clause_prev[8][139] & 1'b1;
			partial_clause[8][140] 	= partial_clause_prev[8][140] & 1'b1;
			partial_clause[8][141] 	= partial_clause_prev[8][141] & 1'b1;
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & 1'b1;
			partial_clause[8][144] 	= partial_clause_prev[8][144] & 1'b1;
			partial_clause[8][145] 	= partial_clause_prev[8][145] & 1'b1;
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & 1'b1;
			partial_clause[8][148] 	= partial_clause_prev[8][148] & 1'b1;
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & 1'b1;
			partial_clause[8][151] 	= partial_clause_prev[8][151] & 1'b1;
			partial_clause[8][152] 	= partial_clause_prev[8][152] & 1'b1;
			partial_clause[8][153] 	= partial_clause_prev[8][153] & 1'b1;
			partial_clause[8][154] 	= partial_clause_prev[8][154] & 1'b1;
			partial_clause[8][155] 	= partial_clause_prev[8][155] & 1'b1;
			partial_clause[8][156] 	= partial_clause_prev[8][156] & 1'b1;
			partial_clause[8][157] 	= partial_clause_prev[8][157] & 1'b1;
			partial_clause[8][158] 	= partial_clause_prev[8][158] & 1'b1;
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & 1'b1;
			partial_clause[8][161] 	= partial_clause_prev[8][161] & 1'b1;
			partial_clause[8][162] 	= partial_clause_prev[8][162] & 1'b1;
			partial_clause[8][163] 	= partial_clause_prev[8][163] & 1'b1;
			partial_clause[8][164] 	= partial_clause_prev[8][164] & 1'b1;
			partial_clause[8][165] 	= partial_clause_prev[8][165] & 1'b1;
			partial_clause[8][166] 	= partial_clause_prev[8][166] & 1'b1;
			partial_clause[8][167] 	= partial_clause_prev[8][167] & 1'b1;
			partial_clause[8][168] 	= partial_clause_prev[8][168] & 1'b1;
			partial_clause[8][169] 	= partial_clause_prev[8][169] & 1'b1;
			partial_clause[8][170] 	= partial_clause_prev[8][170] & 1'b1;
			partial_clause[8][171] 	= partial_clause_prev[8][171] & 1'b1;
			partial_clause[8][172] 	= partial_clause_prev[8][172] & 1'b1;
			partial_clause[8][173] 	= partial_clause_prev[8][173] & 1'b1;
			partial_clause[8][174] 	= partial_clause_prev[8][174] & 1'b1;
			partial_clause[8][175] 	= partial_clause_prev[8][175] & 1'b1;
			partial_clause[8][176] 	= partial_clause_prev[8][176] & 1'b1;
			partial_clause[8][177] 	= partial_clause_prev[8][177] & 1'b1;
			partial_clause[8][178] 	= partial_clause_prev[8][178] & 1'b1;
			partial_clause[8][179] 	= partial_clause_prev[8][179] & 1'b1;
			partial_clause[8][180] 	= partial_clause_prev[8][180] & x[60];
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & ~x[53];
			partial_clause[8][183] 	= partial_clause_prev[8][183] & ~x[6];
			partial_clause[8][184] 	= partial_clause_prev[8][184] & 1'b1;
			partial_clause[8][185] 	= partial_clause_prev[8][185] & 1'b1;
			partial_clause[8][186] 	= partial_clause_prev[8][186] & 1'b1;
			partial_clause[8][187] 	= partial_clause_prev[8][187] & x[4];
			partial_clause[8][188] 	= partial_clause_prev[8][188] & 1'b1;
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & 1'b1;
			partial_clause[8][191] 	= partial_clause_prev[8][191] & 1'b1;
			partial_clause[8][192] 	= partial_clause_prev[8][192] & 1'b1;
			partial_clause[8][193] 	= partial_clause_prev[8][193] & 1'b1;
			partial_clause[8][194] 	= partial_clause_prev[8][194] & 1'b1;
			partial_clause[8][195] 	= partial_clause_prev[8][195] & 1'b1;
			partial_clause[8][196] 	= partial_clause_prev[8][196] & 1'b1;
			partial_clause[8][197] 	= partial_clause_prev[8][197] & 1'b1;
			partial_clause[8][198] 	= partial_clause_prev[8][198] & 1'b1;
			partial_clause[8][199] 	= partial_clause_prev[8][199] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & x[3];
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & x[60];
			partial_clause[9][18] 	= partial_clause_prev[9][18] & x[19] & ~x[40] & ~x[41];
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & ~x[41];
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & ~x[29];
			partial_clause[9][30] 	= partial_clause_prev[9][30] & x[18];
			partial_clause[9][31] 	= partial_clause_prev[9][31] & x[17] & ~x[26];
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & ~x[40];
			partial_clause[9][35] 	= partial_clause_prev[9][35] & x[17];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & x[17];
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & ~x[13] & ~x[39];
			partial_clause[9][49] 	= partial_clause_prev[9][49] & x[20] & ~x[41];
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & x[20];
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & ~x[14] & x[19];
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & x[20];
			partial_clause[9][66] 	= partial_clause_prev[9][66] & x[6];
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & ~x[14] & ~x[15] & x[20];
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & ~x[13] & x[20];
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & x[16];
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & x[47];
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & ~x[13] & ~x[27];
			partial_clause[9][85] 	= partial_clause_prev[9][85] & ~x[13] & x[18];
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & x[32];
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & ~x[13] & x[19] & ~x[40];
			partial_clause[9][100] 	= partial_clause_prev[9][100] & 1'b1;
			partial_clause[9][101] 	= partial_clause_prev[9][101] & ~x[48];
			partial_clause[9][102] 	= partial_clause_prev[9][102] & 1'b1;
			partial_clause[9][103] 	= partial_clause_prev[9][103] & 1'b1;
			partial_clause[9][104] 	= partial_clause_prev[9][104] & 1'b1;
			partial_clause[9][105] 	= partial_clause_prev[9][105] & 1'b1;
			partial_clause[9][106] 	= partial_clause_prev[9][106] & 1'b1;
			partial_clause[9][107] 	= partial_clause_prev[9][107] & 1'b1;
			partial_clause[9][108] 	= partial_clause_prev[9][108] & 1'b1;
			partial_clause[9][109] 	= partial_clause_prev[9][109] & 1'b1;
			partial_clause[9][110] 	= partial_clause_prev[9][110] & 1'b1;
			partial_clause[9][111] 	= partial_clause_prev[9][111] & 1'b1;
			partial_clause[9][112] 	= partial_clause_prev[9][112] & 1'b1;
			partial_clause[9][113] 	= partial_clause_prev[9][113] & ~x[20] & ~x[48];
			partial_clause[9][114] 	= partial_clause_prev[9][114] & 1'b1;
			partial_clause[9][115] 	= partial_clause_prev[9][115] & x[27];
			partial_clause[9][116] 	= partial_clause_prev[9][116] & 1'b1;
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & ~x[20] & ~x[48];
			partial_clause[9][119] 	= partial_clause_prev[9][119] & 1'b1;
			partial_clause[9][120] 	= partial_clause_prev[9][120] & 1'b1;
			partial_clause[9][121] 	= partial_clause_prev[9][121] & 1'b1;
			partial_clause[9][122] 	= partial_clause_prev[9][122] & 1'b1;
			partial_clause[9][123] 	= partial_clause_prev[9][123] & 1'b1;
			partial_clause[9][124] 	= partial_clause_prev[9][124] & 1'b1;
			partial_clause[9][125] 	= partial_clause_prev[9][125] & 1'b1;
			partial_clause[9][126] 	= partial_clause_prev[9][126] & x[1];
			partial_clause[9][127] 	= partial_clause_prev[9][127] & 1'b1;
			partial_clause[9][128] 	= partial_clause_prev[9][128] & 1'b1;
			partial_clause[9][129] 	= partial_clause_prev[9][129] & 1'b1;
			partial_clause[9][130] 	= partial_clause_prev[9][130] & x[27];
			partial_clause[9][131] 	= partial_clause_prev[9][131] & x[11];
			partial_clause[9][132] 	= partial_clause_prev[9][132] & 1'b1;
			partial_clause[9][133] 	= partial_clause_prev[9][133] & 1'b1;
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & 1'b1;
			partial_clause[9][138] 	= partial_clause_prev[9][138] & 1'b1;
			partial_clause[9][139] 	= partial_clause_prev[9][139] & 1'b1;
			partial_clause[9][140] 	= partial_clause_prev[9][140] & x[37];
			partial_clause[9][141] 	= partial_clause_prev[9][141] & 1'b1;
			partial_clause[9][142] 	= partial_clause_prev[9][142] & 1'b1;
			partial_clause[9][143] 	= partial_clause_prev[9][143] & 1'b1;
			partial_clause[9][144] 	= partial_clause_prev[9][144] & ~x[20] & ~x[48];
			partial_clause[9][145] 	= partial_clause_prev[9][145] & 1'b1;
			partial_clause[9][146] 	= partial_clause_prev[9][146] & 1'b1;
			partial_clause[9][147] 	= partial_clause_prev[9][147] & 1'b1;
			partial_clause[9][148] 	= partial_clause_prev[9][148] & 1'b1;
			partial_clause[9][149] 	= partial_clause_prev[9][149] & 1'b1;
			partial_clause[9][150] 	= partial_clause_prev[9][150] & 1'b1;
			partial_clause[9][151] 	= partial_clause_prev[9][151] & 1'b1;
			partial_clause[9][152] 	= partial_clause_prev[9][152] & 1'b1;
			partial_clause[9][153] 	= partial_clause_prev[9][153] & 1'b1;
			partial_clause[9][154] 	= partial_clause_prev[9][154] & 1'b1;
			partial_clause[9][155] 	= partial_clause_prev[9][155] & ~x[19] & ~x[47];
			partial_clause[9][156] 	= partial_clause_prev[9][156] & x[11];
			partial_clause[9][157] 	= partial_clause_prev[9][157] & 1'b1;
			partial_clause[9][158] 	= partial_clause_prev[9][158] & 1'b1;
			partial_clause[9][159] 	= partial_clause_prev[9][159] & 1'b1;
			partial_clause[9][160] 	= partial_clause_prev[9][160] & 1'b1;
			partial_clause[9][161] 	= partial_clause_prev[9][161] & 1'b1;
			partial_clause[9][162] 	= partial_clause_prev[9][162] & x[55];
			partial_clause[9][163] 	= partial_clause_prev[9][163] & 1'b1;
			partial_clause[9][164] 	= partial_clause_prev[9][164] & ~x[19] & ~x[47];
			partial_clause[9][165] 	= partial_clause_prev[9][165] & 1'b1;
			partial_clause[9][166] 	= partial_clause_prev[9][166] & x[26];
			partial_clause[9][167] 	= partial_clause_prev[9][167] & 1'b1;
			partial_clause[9][168] 	= partial_clause_prev[9][168] & 1'b1;
			partial_clause[9][169] 	= partial_clause_prev[9][169] & x[39];
			partial_clause[9][170] 	= partial_clause_prev[9][170] & 1'b1;
			partial_clause[9][171] 	= partial_clause_prev[9][171] & 1'b1;
			partial_clause[9][172] 	= partial_clause_prev[9][172] & 1'b1;
			partial_clause[9][173] 	= partial_clause_prev[9][173] & 1'b1;
			partial_clause[9][174] 	= partial_clause_prev[9][174] & 1'b1;
			partial_clause[9][175] 	= partial_clause_prev[9][175] & ~x[19] & ~x[46];
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & 1'b1;
			partial_clause[9][178] 	= partial_clause_prev[9][178] & 1'b1;
			partial_clause[9][179] 	= partial_clause_prev[9][179] & 1'b1;
			partial_clause[9][180] 	= partial_clause_prev[9][180] & 1'b1;
			partial_clause[9][181] 	= partial_clause_prev[9][181] & 1'b1;
			partial_clause[9][182] 	= partial_clause_prev[9][182] & 1'b1;
			partial_clause[9][183] 	= partial_clause_prev[9][183] & 1'b1;
			partial_clause[9][184] 	= partial_clause_prev[9][184] & 1'b1;
			partial_clause[9][185] 	= partial_clause_prev[9][185] & 1'b1;
			partial_clause[9][186] 	= partial_clause_prev[9][186] & 1'b1;
			partial_clause[9][187] 	= partial_clause_prev[9][187] & ~x[19];
			partial_clause[9][188] 	= partial_clause_prev[9][188] & 1'b1;
			partial_clause[9][189] 	= partial_clause_prev[9][189] & 1'b1;
			partial_clause[9][190] 	= partial_clause_prev[9][190] & 1'b1;
			partial_clause[9][191] 	= partial_clause_prev[9][191] & 1'b1;
			partial_clause[9][192] 	= partial_clause_prev[9][192] & 1'b1;
			partial_clause[9][193] 	= partial_clause_prev[9][193] & 1'b1;
			partial_clause[9][194] 	= partial_clause_prev[9][194] & 1'b1;
			partial_clause[9][195] 	= partial_clause_prev[9][195] & 1'b1;
			partial_clause[9][196] 	= partial_clause_prev[9][196] & 1'b1;
			partial_clause[9][197] 	= partial_clause_prev[9][197] & 1'b1;
			partial_clause[9][198] 	= partial_clause_prev[9][198] & 1'b1;
			partial_clause[9][199] 	= partial_clause_prev[9][199] & 1'b1;
		end
	end
endmodule


module HCB_4 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & x[15];
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & ~x[37];
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & ~x[2];
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & ~x[38];
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & ~x[60];
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & x[13];
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & ~x[57];
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & x[42];
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & ~x[3] & x[44];
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & x[46];
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & x[16];
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & ~x[52];
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & ~x[39];
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & x[12];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & ~x[46];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			partial_clause[0][100] 	= partial_clause_prev[0][100] & 1'b1;
			partial_clause[0][101] 	= partial_clause_prev[0][101] & 1'b1;
			partial_clause[0][102] 	= partial_clause_prev[0][102] & 1'b1;
			partial_clause[0][103] 	= partial_clause_prev[0][103] & 1'b1;
			partial_clause[0][104] 	= partial_clause_prev[0][104] & ~x[42] & ~x[43];
			partial_clause[0][105] 	= partial_clause_prev[0][105] & 1'b1;
			partial_clause[0][106] 	= partial_clause_prev[0][106] & 1'b1;
			partial_clause[0][107] 	= partial_clause_prev[0][107] & 1'b1;
			partial_clause[0][108] 	= partial_clause_prev[0][108] & 1'b1;
			partial_clause[0][109] 	= partial_clause_prev[0][109] & 1'b1;
			partial_clause[0][110] 	= partial_clause_prev[0][110] & 1'b1;
			partial_clause[0][111] 	= partial_clause_prev[0][111] & ~x[38];
			partial_clause[0][112] 	= partial_clause_prev[0][112] & 1'b1;
			partial_clause[0][113] 	= partial_clause_prev[0][113] & 1'b1;
			partial_clause[0][114] 	= partial_clause_prev[0][114] & 1'b1;
			partial_clause[0][115] 	= partial_clause_prev[0][115] & 1'b1;
			partial_clause[0][116] 	= partial_clause_prev[0][116] & ~x[12];
			partial_clause[0][117] 	= partial_clause_prev[0][117] & 1'b1;
			partial_clause[0][118] 	= partial_clause_prev[0][118] & 1'b1;
			partial_clause[0][119] 	= partial_clause_prev[0][119] & ~x[38] & ~x[63];
			partial_clause[0][120] 	= partial_clause_prev[0][120] & 1'b1;
			partial_clause[0][121] 	= partial_clause_prev[0][121] & 1'b1;
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & 1'b1;
			partial_clause[0][124] 	= partial_clause_prev[0][124] & 1'b1;
			partial_clause[0][125] 	= partial_clause_prev[0][125] & ~x[16] & ~x[42];
			partial_clause[0][126] 	= partial_clause_prev[0][126] & 1'b1;
			partial_clause[0][127] 	= partial_clause_prev[0][127] & ~x[10] & ~x[17];
			partial_clause[0][128] 	= partial_clause_prev[0][128] & 1'b1;
			partial_clause[0][129] 	= partial_clause_prev[0][129] & 1'b1;
			partial_clause[0][130] 	= partial_clause_prev[0][130] & 1'b1;
			partial_clause[0][131] 	= partial_clause_prev[0][131] & 1'b1;
			partial_clause[0][132] 	= partial_clause_prev[0][132] & 1'b1;
			partial_clause[0][133] 	= partial_clause_prev[0][133] & 1'b1;
			partial_clause[0][134] 	= partial_clause_prev[0][134] & 1'b1;
			partial_clause[0][135] 	= partial_clause_prev[0][135] & 1'b1;
			partial_clause[0][136] 	= partial_clause_prev[0][136] & 1'b1;
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & 1'b1;
			partial_clause[0][139] 	= partial_clause_prev[0][139] & ~x[9];
			partial_clause[0][140] 	= partial_clause_prev[0][140] & 1'b1;
			partial_clause[0][141] 	= partial_clause_prev[0][141] & ~x[12] & ~x[13];
			partial_clause[0][142] 	= partial_clause_prev[0][142] & 1'b1;
			partial_clause[0][143] 	= partial_clause_prev[0][143] & 1'b1;
			partial_clause[0][144] 	= partial_clause_prev[0][144] & 1'b1;
			partial_clause[0][145] 	= partial_clause_prev[0][145] & 1'b1;
			partial_clause[0][146] 	= partial_clause_prev[0][146] & 1'b1;
			partial_clause[0][147] 	= partial_clause_prev[0][147] & 1'b1;
			partial_clause[0][148] 	= partial_clause_prev[0][148] & 1'b1;
			partial_clause[0][149] 	= partial_clause_prev[0][149] & 1'b1;
			partial_clause[0][150] 	= partial_clause_prev[0][150] & 1'b1;
			partial_clause[0][151] 	= partial_clause_prev[0][151] & 1'b1;
			partial_clause[0][152] 	= partial_clause_prev[0][152] & ~x[12] & ~x[14];
			partial_clause[0][153] 	= partial_clause_prev[0][153] & 1'b1;
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & ~x[37];
			partial_clause[0][156] 	= partial_clause_prev[0][156] & ~x[11];
			partial_clause[0][157] 	= partial_clause_prev[0][157] & 1'b1;
			partial_clause[0][158] 	= partial_clause_prev[0][158] & ~x[37];
			partial_clause[0][159] 	= partial_clause_prev[0][159] & ~x[41];
			partial_clause[0][160] 	= partial_clause_prev[0][160] & 1'b1;
			partial_clause[0][161] 	= partial_clause_prev[0][161] & ~x[14];
			partial_clause[0][162] 	= partial_clause_prev[0][162] & 1'b1;
			partial_clause[0][163] 	= partial_clause_prev[0][163] & 1'b1;
			partial_clause[0][164] 	= partial_clause_prev[0][164] & 1'b1;
			partial_clause[0][165] 	= partial_clause_prev[0][165] & 1'b1;
			partial_clause[0][166] 	= partial_clause_prev[0][166] & 1'b1;
			partial_clause[0][167] 	= partial_clause_prev[0][167] & 1'b1;
			partial_clause[0][168] 	= partial_clause_prev[0][168] & x[50];
			partial_clause[0][169] 	= partial_clause_prev[0][169] & 1'b1;
			partial_clause[0][170] 	= partial_clause_prev[0][170] & 1'b1;
			partial_clause[0][171] 	= partial_clause_prev[0][171] & 1'b1;
			partial_clause[0][172] 	= partial_clause_prev[0][172] & 1'b1;
			partial_clause[0][173] 	= partial_clause_prev[0][173] & ~x[38];
			partial_clause[0][174] 	= partial_clause_prev[0][174] & 1'b1;
			partial_clause[0][175] 	= partial_clause_prev[0][175] & 1'b1;
			partial_clause[0][176] 	= partial_clause_prev[0][176] & 1'b1;
			partial_clause[0][177] 	= partial_clause_prev[0][177] & ~x[63];
			partial_clause[0][178] 	= partial_clause_prev[0][178] & 1'b1;
			partial_clause[0][179] 	= partial_clause_prev[0][179] & 1'b1;
			partial_clause[0][180] 	= partial_clause_prev[0][180] & 1'b1;
			partial_clause[0][181] 	= partial_clause_prev[0][181] & 1'b1;
			partial_clause[0][182] 	= partial_clause_prev[0][182] & 1'b1;
			partial_clause[0][183] 	= partial_clause_prev[0][183] & 1'b1;
			partial_clause[0][184] 	= partial_clause_prev[0][184] & 1'b1;
			partial_clause[0][185] 	= partial_clause_prev[0][185] & 1'b1;
			partial_clause[0][186] 	= partial_clause_prev[0][186] & 1'b1;
			partial_clause[0][187] 	= partial_clause_prev[0][187] & ~x[41];
			partial_clause[0][188] 	= partial_clause_prev[0][188] & 1'b1;
			partial_clause[0][189] 	= partial_clause_prev[0][189] & 1'b1;
			partial_clause[0][190] 	= partial_clause_prev[0][190] & 1'b1;
			partial_clause[0][191] 	= partial_clause_prev[0][191] & 1'b1;
			partial_clause[0][192] 	= partial_clause_prev[0][192] & 1'b1;
			partial_clause[0][193] 	= partial_clause_prev[0][193] & ~x[41];
			partial_clause[0][194] 	= partial_clause_prev[0][194] & 1'b1;
			partial_clause[0][195] 	= partial_clause_prev[0][195] & 1'b1;
			partial_clause[0][196] 	= partial_clause_prev[0][196] & 1'b1;
			partial_clause[0][197] 	= partial_clause_prev[0][197] & 1'b1;
			partial_clause[0][198] 	= partial_clause_prev[0][198] & ~x[17] & ~x[18] & ~x[26] & ~x[41] & ~x[43];
			partial_clause[0][199] 	= partial_clause_prev[0][199] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & ~x[36];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & ~x[14];
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & ~x[42];
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & ~x[42];
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & ~x[13];
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & ~x[42];
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & x[37];
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & ~x[41];
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & ~x[7];
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & x[13];
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & ~x[13];
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & 1'b1;
			partial_clause[1][59] 	= partial_clause_prev[1][59] & ~x[46];
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & ~x[7] & x[40];
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & x[40];
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & ~x[16] & x[38] & ~x[57];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & ~x[13] & ~x[42];
			partial_clause[1][78] 	= partial_clause_prev[1][78] & ~x[9];
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & ~x[17];
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & ~x[14] & ~x[42];
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & x[37];
			partial_clause[1][90] 	= partial_clause_prev[1][90] & ~x[20];
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & ~x[36];
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			partial_clause[1][100] 	= partial_clause_prev[1][100] & 1'b1;
			partial_clause[1][101] 	= partial_clause_prev[1][101] & ~x[11];
			partial_clause[1][102] 	= partial_clause_prev[1][102] & 1'b1;
			partial_clause[1][103] 	= partial_clause_prev[1][103] & 1'b1;
			partial_clause[1][104] 	= partial_clause_prev[1][104] & 1'b1;
			partial_clause[1][105] 	= partial_clause_prev[1][105] & 1'b1;
			partial_clause[1][106] 	= partial_clause_prev[1][106] & 1'b1;
			partial_clause[1][107] 	= partial_clause_prev[1][107] & 1'b1;
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & ~x[38];
			partial_clause[1][110] 	= partial_clause_prev[1][110] & 1'b1;
			partial_clause[1][111] 	= partial_clause_prev[1][111] & 1'b1;
			partial_clause[1][112] 	= partial_clause_prev[1][112] & 1'b1;
			partial_clause[1][113] 	= partial_clause_prev[1][113] & 1'b1;
			partial_clause[1][114] 	= partial_clause_prev[1][114] & 1'b1;
			partial_clause[1][115] 	= partial_clause_prev[1][115] & 1'b1;
			partial_clause[1][116] 	= partial_clause_prev[1][116] & 1'b1;
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & ~x[39];
			partial_clause[1][119] 	= partial_clause_prev[1][119] & x[59];
			partial_clause[1][120] 	= partial_clause_prev[1][120] & 1'b1;
			partial_clause[1][121] 	= partial_clause_prev[1][121] & 1'b1;
			partial_clause[1][122] 	= partial_clause_prev[1][122] & x[34];
			partial_clause[1][123] 	= partial_clause_prev[1][123] & 1'b1;
			partial_clause[1][124] 	= partial_clause_prev[1][124] & ~x[9];
			partial_clause[1][125] 	= partial_clause_prev[1][125] & 1'b1;
			partial_clause[1][126] 	= partial_clause_prev[1][126] & 1'b1;
			partial_clause[1][127] 	= partial_clause_prev[1][127] & 1'b1;
			partial_clause[1][128] 	= partial_clause_prev[1][128] & 1'b1;
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & x[42];
			partial_clause[1][131] 	= partial_clause_prev[1][131] & 1'b1;
			partial_clause[1][132] 	= partial_clause_prev[1][132] & 1'b1;
			partial_clause[1][133] 	= partial_clause_prev[1][133] & 1'b1;
			partial_clause[1][134] 	= partial_clause_prev[1][134] & 1'b1;
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & 1'b1;
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & x[34];
			partial_clause[1][139] 	= partial_clause_prev[1][139] & 1'b1;
			partial_clause[1][140] 	= partial_clause_prev[1][140] & 1'b1;
			partial_clause[1][141] 	= partial_clause_prev[1][141] & 1'b1;
			partial_clause[1][142] 	= partial_clause_prev[1][142] & 1'b1;
			partial_clause[1][143] 	= partial_clause_prev[1][143] & 1'b1;
			partial_clause[1][144] 	= partial_clause_prev[1][144] & 1'b1;
			partial_clause[1][145] 	= partial_clause_prev[1][145] & 1'b1;
			partial_clause[1][146] 	= partial_clause_prev[1][146] & ~x[9];
			partial_clause[1][147] 	= partial_clause_prev[1][147] & ~x[36];
			partial_clause[1][148] 	= partial_clause_prev[1][148] & 1'b1;
			partial_clause[1][149] 	= partial_clause_prev[1][149] & 1'b1;
			partial_clause[1][150] 	= partial_clause_prev[1][150] & 1'b1;
			partial_clause[1][151] 	= partial_clause_prev[1][151] & 1'b1;
			partial_clause[1][152] 	= partial_clause_prev[1][152] & 1'b1;
			partial_clause[1][153] 	= partial_clause_prev[1][153] & 1'b1;
			partial_clause[1][154] 	= partial_clause_prev[1][154] & 1'b1;
			partial_clause[1][155] 	= partial_clause_prev[1][155] & 1'b1;
			partial_clause[1][156] 	= partial_clause_prev[1][156] & 1'b1;
			partial_clause[1][157] 	= partial_clause_prev[1][157] & 1'b1;
			partial_clause[1][158] 	= partial_clause_prev[1][158] & 1'b1;
			partial_clause[1][159] 	= partial_clause_prev[1][159] & 1'b1;
			partial_clause[1][160] 	= partial_clause_prev[1][160] & 1'b1;
			partial_clause[1][161] 	= partial_clause_prev[1][161] & 1'b1;
			partial_clause[1][162] 	= partial_clause_prev[1][162] & 1'b1;
			partial_clause[1][163] 	= partial_clause_prev[1][163] & 1'b1;
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & 1'b1;
			partial_clause[1][166] 	= partial_clause_prev[1][166] & 1'b1;
			partial_clause[1][167] 	= partial_clause_prev[1][167] & 1'b1;
			partial_clause[1][168] 	= partial_clause_prev[1][168] & 1'b1;
			partial_clause[1][169] 	= partial_clause_prev[1][169] & 1'b1;
			partial_clause[1][170] 	= partial_clause_prev[1][170] & 1'b1;
			partial_clause[1][171] 	= partial_clause_prev[1][171] & 1'b1;
			partial_clause[1][172] 	= partial_clause_prev[1][172] & x[61];
			partial_clause[1][173] 	= partial_clause_prev[1][173] & ~x[38] & x[63];
			partial_clause[1][174] 	= partial_clause_prev[1][174] & x[45];
			partial_clause[1][175] 	= partial_clause_prev[1][175] & ~x[39];
			partial_clause[1][176] 	= partial_clause_prev[1][176] & 1'b1;
			partial_clause[1][177] 	= partial_clause_prev[1][177] & 1'b1;
			partial_clause[1][178] 	= partial_clause_prev[1][178] & 1'b1;
			partial_clause[1][179] 	= partial_clause_prev[1][179] & 1'b1;
			partial_clause[1][180] 	= partial_clause_prev[1][180] & ~x[36];
			partial_clause[1][181] 	= partial_clause_prev[1][181] & 1'b1;
			partial_clause[1][182] 	= partial_clause_prev[1][182] & 1'b1;
			partial_clause[1][183] 	= partial_clause_prev[1][183] & 1'b1;
			partial_clause[1][184] 	= partial_clause_prev[1][184] & 1'b1;
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & 1'b1;
			partial_clause[1][187] 	= partial_clause_prev[1][187] & 1'b1;
			partial_clause[1][188] 	= partial_clause_prev[1][188] & ~x[8];
			partial_clause[1][189] 	= partial_clause_prev[1][189] & 1'b1;
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & 1'b1;
			partial_clause[1][192] 	= partial_clause_prev[1][192] & 1'b1;
			partial_clause[1][193] 	= partial_clause_prev[1][193] & ~x[39];
			partial_clause[1][194] 	= partial_clause_prev[1][194] & 1'b1;
			partial_clause[1][195] 	= partial_clause_prev[1][195] & 1'b1;
			partial_clause[1][196] 	= partial_clause_prev[1][196] & ~x[38];
			partial_clause[1][197] 	= partial_clause_prev[1][197] & 1'b1;
			partial_clause[1][198] 	= partial_clause_prev[1][198] & ~x[9];
			partial_clause[1][199] 	= partial_clause_prev[1][199] & ~x[38];
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & ~x[5] & ~x[34] & ~x[35] & ~x[61];
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & ~x[61];
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & ~x[5] & ~x[32] & ~x[57] & ~x[63];
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & ~x[2] & ~x[34];
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & ~x[7] & ~x[59] & ~x[61];
			partial_clause[2][35] 	= partial_clause_prev[2][35] & ~x[38];
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & ~x[9] & ~x[36] & ~x[38] & ~x[61] & ~x[62];
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & ~x[6] & ~x[7];
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & 1'b1;
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & ~x[36] & ~x[60];
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & ~x[61] & ~x[62];
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & ~x[6] & ~x[31] & ~x[58];
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & ~x[62];
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			partial_clause[2][100] 	= partial_clause_prev[2][100] & 1'b1;
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & 1'b1;
			partial_clause[2][103] 	= partial_clause_prev[2][103] & 1'b1;
			partial_clause[2][104] 	= partial_clause_prev[2][104] & 1'b1;
			partial_clause[2][105] 	= partial_clause_prev[2][105] & ~x[33] & x[37];
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & 1'b1;
			partial_clause[2][108] 	= partial_clause_prev[2][108] & x[31];
			partial_clause[2][109] 	= partial_clause_prev[2][109] & 1'b1;
			partial_clause[2][110] 	= partial_clause_prev[2][110] & x[59];
			partial_clause[2][111] 	= partial_clause_prev[2][111] & 1'b1;
			partial_clause[2][112] 	= partial_clause_prev[2][112] & x[63];
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & 1'b1;
			partial_clause[2][115] 	= partial_clause_prev[2][115] & 1'b1;
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & x[59];
			partial_clause[2][118] 	= partial_clause_prev[2][118] & 1'b1;
			partial_clause[2][119] 	= partial_clause_prev[2][119] & x[61];
			partial_clause[2][120] 	= partial_clause_prev[2][120] & x[63];
			partial_clause[2][121] 	= partial_clause_prev[2][121] & 1'b1;
			partial_clause[2][122] 	= partial_clause_prev[2][122] & 1'b1;
			partial_clause[2][123] 	= partial_clause_prev[2][123] & 1'b1;
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & 1'b1;
			partial_clause[2][126] 	= partial_clause_prev[2][126] & 1'b1;
			partial_clause[2][127] 	= partial_clause_prev[2][127] & x[61];
			partial_clause[2][128] 	= partial_clause_prev[2][128] & x[36];
			partial_clause[2][129] 	= partial_clause_prev[2][129] & 1'b1;
			partial_clause[2][130] 	= partial_clause_prev[2][130] & 1'b1;
			partial_clause[2][131] 	= partial_clause_prev[2][131] & 1'b1;
			partial_clause[2][132] 	= partial_clause_prev[2][132] & x[61];
			partial_clause[2][133] 	= partial_clause_prev[2][133] & 1'b1;
			partial_clause[2][134] 	= partial_clause_prev[2][134] & 1'b1;
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & 1'b1;
			partial_clause[2][137] 	= partial_clause_prev[2][137] & 1'b1;
			partial_clause[2][138] 	= partial_clause_prev[2][138] & 1'b1;
			partial_clause[2][139] 	= partial_clause_prev[2][139] & 1'b1;
			partial_clause[2][140] 	= partial_clause_prev[2][140] & 1'b1;
			partial_clause[2][141] 	= partial_clause_prev[2][141] & 1'b1;
			partial_clause[2][142] 	= partial_clause_prev[2][142] & x[59];
			partial_clause[2][143] 	= partial_clause_prev[2][143] & 1'b1;
			partial_clause[2][144] 	= partial_clause_prev[2][144] & 1'b1;
			partial_clause[2][145] 	= partial_clause_prev[2][145] & 1'b1;
			partial_clause[2][146] 	= partial_clause_prev[2][146] & 1'b1;
			partial_clause[2][147] 	= partial_clause_prev[2][147] & 1'b1;
			partial_clause[2][148] 	= partial_clause_prev[2][148] & 1'b1;
			partial_clause[2][149] 	= partial_clause_prev[2][149] & 1'b1;
			partial_clause[2][150] 	= partial_clause_prev[2][150] & 1'b1;
			partial_clause[2][151] 	= partial_clause_prev[2][151] & 1'b1;
			partial_clause[2][152] 	= partial_clause_prev[2][152] & 1'b1;
			partial_clause[2][153] 	= partial_clause_prev[2][153] & 1'b1;
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & 1'b1;
			partial_clause[2][156] 	= partial_clause_prev[2][156] & 1'b1;
			partial_clause[2][157] 	= partial_clause_prev[2][157] & x[62];
			partial_clause[2][158] 	= partial_clause_prev[2][158] & x[57];
			partial_clause[2][159] 	= partial_clause_prev[2][159] & x[60];
			partial_clause[2][160] 	= partial_clause_prev[2][160] & x[59];
			partial_clause[2][161] 	= partial_clause_prev[2][161] & 1'b1;
			partial_clause[2][162] 	= partial_clause_prev[2][162] & 1'b1;
			partial_clause[2][163] 	= partial_clause_prev[2][163] & 1'b1;
			partial_clause[2][164] 	= partial_clause_prev[2][164] & x[62];
			partial_clause[2][165] 	= partial_clause_prev[2][165] & 1'b1;
			partial_clause[2][166] 	= partial_clause_prev[2][166] & 1'b1;
			partial_clause[2][167] 	= partial_clause_prev[2][167] & 1'b1;
			partial_clause[2][168] 	= partial_clause_prev[2][168] & 1'b1;
			partial_clause[2][169] 	= partial_clause_prev[2][169] & 1'b1;
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & 1'b1;
			partial_clause[2][173] 	= partial_clause_prev[2][173] & 1'b1;
			partial_clause[2][174] 	= partial_clause_prev[2][174] & 1'b1;
			partial_clause[2][175] 	= partial_clause_prev[2][175] & 1'b1;
			partial_clause[2][176] 	= partial_clause_prev[2][176] & 1'b1;
			partial_clause[2][177] 	= partial_clause_prev[2][177] & 1'b1;
			partial_clause[2][178] 	= partial_clause_prev[2][178] & 1'b1;
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & 1'b1;
			partial_clause[2][181] 	= partial_clause_prev[2][181] & 1'b1;
			partial_clause[2][182] 	= partial_clause_prev[2][182] & x[63];
			partial_clause[2][183] 	= partial_clause_prev[2][183] & x[62];
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & 1'b1;
			partial_clause[2][186] 	= partial_clause_prev[2][186] & ~x[33];
			partial_clause[2][187] 	= partial_clause_prev[2][187] & x[21];
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & ~x[33];
			partial_clause[2][190] 	= partial_clause_prev[2][190] & 1'b1;
			partial_clause[2][191] 	= partial_clause_prev[2][191] & 1'b1;
			partial_clause[2][192] 	= partial_clause_prev[2][192] & 1'b1;
			partial_clause[2][193] 	= partial_clause_prev[2][193] & 1'b1;
			partial_clause[2][194] 	= partial_clause_prev[2][194] & 1'b1;
			partial_clause[2][195] 	= partial_clause_prev[2][195] & 1'b1;
			partial_clause[2][196] 	= partial_clause_prev[2][196] & 1'b1;
			partial_clause[2][197] 	= partial_clause_prev[2][197] & 1'b1;
			partial_clause[2][198] 	= partial_clause_prev[2][198] & 1'b1;
			partial_clause[2][199] 	= partial_clause_prev[2][199] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & ~x[63];
			partial_clause[3][1] 	= partial_clause_prev[3][1] & x[9];
			partial_clause[3][2] 	= partial_clause_prev[3][2] & ~x[33];
			partial_clause[3][3] 	= partial_clause_prev[3][3] & ~x[63];
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & ~x[17] & x[38];
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & x[38];
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & x[10];
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & x[13] & ~x[34];
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & ~x[33] & ~x[35];
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & ~x[63];
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & ~x[36] & ~x[62];
			partial_clause[3][38] 	= partial_clause_prev[3][38] & ~x[7] & ~x[30] & ~x[33];
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & ~x[4] & ~x[6] & ~x[8];
			partial_clause[3][41] 	= partial_clause_prev[3][41] & x[13];
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & ~x[7] & ~x[58];
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & ~x[63];
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & x[43];
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & ~x[36];
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & x[11];
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & x[14];
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & 1'b1;
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & ~x[37] & ~x[63];
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & ~x[36] & ~x[62];
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & x[38];
			partial_clause[3][81] 	= partial_clause_prev[3][81] & ~x[5] & ~x[6];
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & x[37];
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & x[39];
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & ~x[62];
			partial_clause[3][96] 	= partial_clause_prev[3][96] & ~x[36];
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & ~x[5] & ~x[6];
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			partial_clause[3][100] 	= partial_clause_prev[3][100] & 1'b1;
			partial_clause[3][101] 	= partial_clause_prev[3][101] & 1'b1;
			partial_clause[3][102] 	= partial_clause_prev[3][102] & 1'b1;
			partial_clause[3][103] 	= partial_clause_prev[3][103] & 1'b1;
			partial_clause[3][104] 	= partial_clause_prev[3][104] & 1'b1;
			partial_clause[3][105] 	= partial_clause_prev[3][105] & x[34] & ~x[37];
			partial_clause[3][106] 	= partial_clause_prev[3][106] & 1'b1;
			partial_clause[3][107] 	= partial_clause_prev[3][107] & 1'b1;
			partial_clause[3][108] 	= partial_clause_prev[3][108] & 1'b1;
			partial_clause[3][109] 	= partial_clause_prev[3][109] & 1'b1;
			partial_clause[3][110] 	= partial_clause_prev[3][110] & 1'b1;
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & 1'b1;
			partial_clause[3][113] 	= partial_clause_prev[3][113] & 1'b1;
			partial_clause[3][114] 	= partial_clause_prev[3][114] & 1'b1;
			partial_clause[3][115] 	= partial_clause_prev[3][115] & 1'b1;
			partial_clause[3][116] 	= partial_clause_prev[3][116] & x[33];
			partial_clause[3][117] 	= partial_clause_prev[3][117] & 1'b1;
			partial_clause[3][118] 	= partial_clause_prev[3][118] & 1'b1;
			partial_clause[3][119] 	= partial_clause_prev[3][119] & 1'b1;
			partial_clause[3][120] 	= partial_clause_prev[3][120] & x[32];
			partial_clause[3][121] 	= partial_clause_prev[3][121] & x[33];
			partial_clause[3][122] 	= partial_clause_prev[3][122] & ~x[38];
			partial_clause[3][123] 	= partial_clause_prev[3][123] & 1'b1;
			partial_clause[3][124] 	= partial_clause_prev[3][124] & 1'b1;
			partial_clause[3][125] 	= partial_clause_prev[3][125] & x[33];
			partial_clause[3][126] 	= partial_clause_prev[3][126] & 1'b1;
			partial_clause[3][127] 	= partial_clause_prev[3][127] & ~x[37];
			partial_clause[3][128] 	= partial_clause_prev[3][128] & ~x[4];
			partial_clause[3][129] 	= partial_clause_prev[3][129] & 1'b1;
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & 1'b1;
			partial_clause[3][132] 	= partial_clause_prev[3][132] & 1'b1;
			partial_clause[3][133] 	= partial_clause_prev[3][133] & 1'b1;
			partial_clause[3][134] 	= partial_clause_prev[3][134] & 1'b1;
			partial_clause[3][135] 	= partial_clause_prev[3][135] & 1'b1;
			partial_clause[3][136] 	= partial_clause_prev[3][136] & 1'b1;
			partial_clause[3][137] 	= partial_clause_prev[3][137] & 1'b1;
			partial_clause[3][138] 	= partial_clause_prev[3][138] & ~x[16];
			partial_clause[3][139] 	= partial_clause_prev[3][139] & 1'b1;
			partial_clause[3][140] 	= partial_clause_prev[3][140] & 1'b1;
			partial_clause[3][141] 	= partial_clause_prev[3][141] & 1'b1;
			partial_clause[3][142] 	= partial_clause_prev[3][142] & 1'b1;
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & 1'b1;
			partial_clause[3][145] 	= partial_clause_prev[3][145] & ~x[5];
			partial_clause[3][146] 	= partial_clause_prev[3][146] & x[60];
			partial_clause[3][147] 	= partial_clause_prev[3][147] & 1'b1;
			partial_clause[3][148] 	= partial_clause_prev[3][148] & 1'b1;
			partial_clause[3][149] 	= partial_clause_prev[3][149] & 1'b1;
			partial_clause[3][150] 	= partial_clause_prev[3][150] & 1'b1;
			partial_clause[3][151] 	= partial_clause_prev[3][151] & ~x[41];
			partial_clause[3][152] 	= partial_clause_prev[3][152] & 1'b1;
			partial_clause[3][153] 	= partial_clause_prev[3][153] & 1'b1;
			partial_clause[3][154] 	= partial_clause_prev[3][154] & 1'b1;
			partial_clause[3][155] 	= partial_clause_prev[3][155] & 1'b1;
			partial_clause[3][156] 	= partial_clause_prev[3][156] & 1'b1;
			partial_clause[3][157] 	= partial_clause_prev[3][157] & 1'b1;
			partial_clause[3][158] 	= partial_clause_prev[3][158] & ~x[40];
			partial_clause[3][159] 	= partial_clause_prev[3][159] & 1'b1;
			partial_clause[3][160] 	= partial_clause_prev[3][160] & 1'b1;
			partial_clause[3][161] 	= partial_clause_prev[3][161] & 1'b1;
			partial_clause[3][162] 	= partial_clause_prev[3][162] & 1'b1;
			partial_clause[3][163] 	= partial_clause_prev[3][163] & 1'b1;
			partial_clause[3][164] 	= partial_clause_prev[3][164] & 1'b1;
			partial_clause[3][165] 	= partial_clause_prev[3][165] & 1'b1;
			partial_clause[3][166] 	= partial_clause_prev[3][166] & 1'b1;
			partial_clause[3][167] 	= partial_clause_prev[3][167] & 1'b1;
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & 1'b1;
			partial_clause[3][170] 	= partial_clause_prev[3][170] & 1'b1;
			partial_clause[3][171] 	= partial_clause_prev[3][171] & 1'b1;
			partial_clause[3][172] 	= partial_clause_prev[3][172] & 1'b1;
			partial_clause[3][173] 	= partial_clause_prev[3][173] & 1'b1;
			partial_clause[3][174] 	= partial_clause_prev[3][174] & 1'b1;
			partial_clause[3][175] 	= partial_clause_prev[3][175] & 1'b1;
			partial_clause[3][176] 	= partial_clause_prev[3][176] & 1'b1;
			partial_clause[3][177] 	= partial_clause_prev[3][177] & x[35];
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & 1'b1;
			partial_clause[3][180] 	= partial_clause_prev[3][180] & x[35];
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & x[60];
			partial_clause[3][183] 	= partial_clause_prev[3][183] & 1'b1;
			partial_clause[3][184] 	= partial_clause_prev[3][184] & 1'b1;
			partial_clause[3][185] 	= partial_clause_prev[3][185] & x[48];
			partial_clause[3][186] 	= partial_clause_prev[3][186] & 1'b1;
			partial_clause[3][187] 	= partial_clause_prev[3][187] & ~x[40];
			partial_clause[3][188] 	= partial_clause_prev[3][188] & 1'b1;
			partial_clause[3][189] 	= partial_clause_prev[3][189] & 1'b1;
			partial_clause[3][190] 	= partial_clause_prev[3][190] & 1'b1;
			partial_clause[3][191] 	= partial_clause_prev[3][191] & 1'b1;
			partial_clause[3][192] 	= partial_clause_prev[3][192] & ~x[9] & x[34];
			partial_clause[3][193] 	= partial_clause_prev[3][193] & 1'b1;
			partial_clause[3][194] 	= partial_clause_prev[3][194] & x[62];
			partial_clause[3][195] 	= partial_clause_prev[3][195] & x[20];
			partial_clause[3][196] 	= partial_clause_prev[3][196] & 1'b1;
			partial_clause[3][197] 	= partial_clause_prev[3][197] & 1'b1;
			partial_clause[3][198] 	= partial_clause_prev[3][198] & 1'b1;
			partial_clause[3][199] 	= partial_clause_prev[3][199] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & ~x[10];
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & ~x[35];
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & ~x[38];
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & ~x[11] & ~x[39];
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[38];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & ~x[33] & x[36];
			partial_clause[4][35] 	= partial_clause_prev[4][35] & ~x[39];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & ~x[12];
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[9];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & ~x[9] & ~x[10];
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & ~x[46];
			partial_clause[4][53] 	= partial_clause_prev[4][53] & ~x[11] & ~x[38];
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & ~x[10];
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & x[63];
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & x[15] & ~x[40];
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & ~x[9];
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & ~x[9] & ~x[38];
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & ~x[11];
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & ~x[38];
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & x[43];
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			partial_clause[4][100] 	= partial_clause_prev[4][100] & 1'b1;
			partial_clause[4][101] 	= partial_clause_prev[4][101] & 1'b1;
			partial_clause[4][102] 	= partial_clause_prev[4][102] & 1'b1;
			partial_clause[4][103] 	= partial_clause_prev[4][103] & 1'b1;
			partial_clause[4][104] 	= partial_clause_prev[4][104] & 1'b1;
			partial_clause[4][105] 	= partial_clause_prev[4][105] & 1'b1;
			partial_clause[4][106] 	= partial_clause_prev[4][106] & 1'b1;
			partial_clause[4][107] 	= partial_clause_prev[4][107] & 1'b1;
			partial_clause[4][108] 	= partial_clause_prev[4][108] & 1'b1;
			partial_clause[4][109] 	= partial_clause_prev[4][109] & 1'b1;
			partial_clause[4][110] 	= partial_clause_prev[4][110] & 1'b1;
			partial_clause[4][111] 	= partial_clause_prev[4][111] & 1'b1;
			partial_clause[4][112] 	= partial_clause_prev[4][112] & 1'b1;
			partial_clause[4][113] 	= partial_clause_prev[4][113] & ~x[41] & ~x[46];
			partial_clause[4][114] 	= partial_clause_prev[4][114] & 1'b1;
			partial_clause[4][115] 	= partial_clause_prev[4][115] & 1'b1;
			partial_clause[4][116] 	= partial_clause_prev[4][116] & ~x[14];
			partial_clause[4][117] 	= partial_clause_prev[4][117] & 1'b1;
			partial_clause[4][118] 	= partial_clause_prev[4][118] & 1'b1;
			partial_clause[4][119] 	= partial_clause_prev[4][119] & 1'b1;
			partial_clause[4][120] 	= partial_clause_prev[4][120] & 1'b1;
			partial_clause[4][121] 	= partial_clause_prev[4][121] & 1'b1;
			partial_clause[4][122] 	= partial_clause_prev[4][122] & ~x[37];
			partial_clause[4][123] 	= partial_clause_prev[4][123] & 1'b1;
			partial_clause[4][124] 	= partial_clause_prev[4][124] & 1'b1;
			partial_clause[4][125] 	= partial_clause_prev[4][125] & 1'b1;
			partial_clause[4][126] 	= partial_clause_prev[4][126] & 1'b1;
			partial_clause[4][127] 	= partial_clause_prev[4][127] & 1'b1;
			partial_clause[4][128] 	= partial_clause_prev[4][128] & 1'b1;
			partial_clause[4][129] 	= partial_clause_prev[4][129] & 1'b1;
			partial_clause[4][130] 	= partial_clause_prev[4][130] & 1'b1;
			partial_clause[4][131] 	= partial_clause_prev[4][131] & 1'b1;
			partial_clause[4][132] 	= partial_clause_prev[4][132] & 1'b1;
			partial_clause[4][133] 	= partial_clause_prev[4][133] & 1'b1;
			partial_clause[4][134] 	= partial_clause_prev[4][134] & 1'b1;
			partial_clause[4][135] 	= partial_clause_prev[4][135] & 1'b1;
			partial_clause[4][136] 	= partial_clause_prev[4][136] & 1'b1;
			partial_clause[4][137] 	= partial_clause_prev[4][137] & 1'b1;
			partial_clause[4][138] 	= partial_clause_prev[4][138] & 1'b1;
			partial_clause[4][139] 	= partial_clause_prev[4][139] & 1'b1;
			partial_clause[4][140] 	= partial_clause_prev[4][140] & 1'b1;
			partial_clause[4][141] 	= partial_clause_prev[4][141] & 1'b1;
			partial_clause[4][142] 	= partial_clause_prev[4][142] & 1'b1;
			partial_clause[4][143] 	= partial_clause_prev[4][143] & x[12] & x[43];
			partial_clause[4][144] 	= partial_clause_prev[4][144] & 1'b1;
			partial_clause[4][145] 	= partial_clause_prev[4][145] & 1'b1;
			partial_clause[4][146] 	= partial_clause_prev[4][146] & 1'b1;
			partial_clause[4][147] 	= partial_clause_prev[4][147] & 1'b1;
			partial_clause[4][148] 	= partial_clause_prev[4][148] & 1'b1;
			partial_clause[4][149] 	= partial_clause_prev[4][149] & 1'b1;
			partial_clause[4][150] 	= partial_clause_prev[4][150] & 1'b1;
			partial_clause[4][151] 	= partial_clause_prev[4][151] & 1'b1;
			partial_clause[4][152] 	= partial_clause_prev[4][152] & 1'b1;
			partial_clause[4][153] 	= partial_clause_prev[4][153] & ~x[45];
			partial_clause[4][154] 	= partial_clause_prev[4][154] & 1'b1;
			partial_clause[4][155] 	= partial_clause_prev[4][155] & ~x[40];
			partial_clause[4][156] 	= partial_clause_prev[4][156] & 1'b1;
			partial_clause[4][157] 	= partial_clause_prev[4][157] & 1'b1;
			partial_clause[4][158] 	= partial_clause_prev[4][158] & 1'b1;
			partial_clause[4][159] 	= partial_clause_prev[4][159] & 1'b1;
			partial_clause[4][160] 	= partial_clause_prev[4][160] & 1'b1;
			partial_clause[4][161] 	= partial_clause_prev[4][161] & 1'b1;
			partial_clause[4][162] 	= partial_clause_prev[4][162] & 1'b1;
			partial_clause[4][163] 	= partial_clause_prev[4][163] & 1'b1;
			partial_clause[4][164] 	= partial_clause_prev[4][164] & 1'b1;
			partial_clause[4][165] 	= partial_clause_prev[4][165] & 1'b1;
			partial_clause[4][166] 	= partial_clause_prev[4][166] & 1'b1;
			partial_clause[4][167] 	= partial_clause_prev[4][167] & 1'b1;
			partial_clause[4][168] 	= partial_clause_prev[4][168] & 1'b1;
			partial_clause[4][169] 	= partial_clause_prev[4][169] & 1'b1;
			partial_clause[4][170] 	= partial_clause_prev[4][170] & 1'b1;
			partial_clause[4][171] 	= partial_clause_prev[4][171] & 1'b1;
			partial_clause[4][172] 	= partial_clause_prev[4][172] & 1'b1;
			partial_clause[4][173] 	= partial_clause_prev[4][173] & 1'b1;
			partial_clause[4][174] 	= partial_clause_prev[4][174] & ~x[36];
			partial_clause[4][175] 	= partial_clause_prev[4][175] & 1'b1;
			partial_clause[4][176] 	= partial_clause_prev[4][176] & 1'b1;
			partial_clause[4][177] 	= partial_clause_prev[4][177] & 1'b1;
			partial_clause[4][178] 	= partial_clause_prev[4][178] & 1'b1;
			partial_clause[4][179] 	= partial_clause_prev[4][179] & 1'b1;
			partial_clause[4][180] 	= partial_clause_prev[4][180] & 1'b1;
			partial_clause[4][181] 	= partial_clause_prev[4][181] & ~x[9] & ~x[36];
			partial_clause[4][182] 	= partial_clause_prev[4][182] & 1'b1;
			partial_clause[4][183] 	= partial_clause_prev[4][183] & x[7] & x[10];
			partial_clause[4][184] 	= partial_clause_prev[4][184] & 1'b1;
			partial_clause[4][185] 	= partial_clause_prev[4][185] & 1'b1;
			partial_clause[4][186] 	= partial_clause_prev[4][186] & 1'b1;
			partial_clause[4][187] 	= partial_clause_prev[4][187] & ~x[63];
			partial_clause[4][188] 	= partial_clause_prev[4][188] & 1'b1;
			partial_clause[4][189] 	= partial_clause_prev[4][189] & 1'b1;
			partial_clause[4][190] 	= partial_clause_prev[4][190] & ~x[62];
			partial_clause[4][191] 	= partial_clause_prev[4][191] & 1'b1;
			partial_clause[4][192] 	= partial_clause_prev[4][192] & 1'b1;
			partial_clause[4][193] 	= partial_clause_prev[4][193] & 1'b1;
			partial_clause[4][194] 	= partial_clause_prev[4][194] & 1'b1;
			partial_clause[4][195] 	= partial_clause_prev[4][195] & x[8];
			partial_clause[4][196] 	= partial_clause_prev[4][196] & 1'b1;
			partial_clause[4][197] 	= partial_clause_prev[4][197] & 1'b1;
			partial_clause[4][198] 	= partial_clause_prev[4][198] & ~x[12] & ~x[14];
			partial_clause[4][199] 	= partial_clause_prev[4][199] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & ~x[42] & ~x[43] & ~x[44] & ~x[46];
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & x[49];
			partial_clause[5][3] 	= partial_clause_prev[5][3] & x[33] & ~x[44] & ~x[46];
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & x[40] & x[42];
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & ~x[12] & ~x[14] & ~x[15] & ~x[17];
			partial_clause[5][12] 	= partial_clause_prev[5][12] & ~x[40] & ~x[42] & ~x[43];
			partial_clause[5][13] 	= partial_clause_prev[5][13] & x[20];
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & x[49];
			partial_clause[5][16] 	= partial_clause_prev[5][16] & x[13] & x[17];
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & x[48];
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & ~x[10] & ~x[11] & ~x[14] & ~x[18];
			partial_clause[5][21] 	= partial_clause_prev[5][21] & x[15];
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & x[36];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & x[49];
			partial_clause[5][26] 	= partial_clause_prev[5][26] & x[20];
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & x[48];
			partial_clause[5][32] 	= partial_clause_prev[5][32] & x[58];
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & ~x[39] & ~x[41] & ~x[44] & ~x[46];
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & ~x[39] & ~x[41] & ~x[43] & ~x[44] & ~x[47];
			partial_clause[5][40] 	= partial_clause_prev[5][40] & ~x[13] & ~x[44];
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & ~x[38] & ~x[41] & ~x[43] & ~x[46];
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & ~x[38] & ~x[40] & ~x[41] & ~x[43];
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & x[50];
			partial_clause[5][49] 	= partial_clause_prev[5][49] & x[49];
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & x[48];
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & ~x[10] & ~x[14] & ~x[17];
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & ~x[42] & ~x[44] & ~x[46] & ~x[47];
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & x[40] & x[41];
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & ~x[41] & ~x[43];
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & x[49];
			partial_clause[5][65] 	= partial_clause_prev[5][65] & ~x[43];
			partial_clause[5][66] 	= partial_clause_prev[5][66] & x[20];
			partial_clause[5][67] 	= partial_clause_prev[5][67] & x[15];
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & ~x[1];
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & x[60];
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & x[49];
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & x[49];
			partial_clause[5][80] 	= partial_clause_prev[5][80] & x[19];
			partial_clause[5][81] 	= partial_clause_prev[5][81] & ~x[10] & ~x[12];
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & x[17] & x[20];
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & ~x[15] & ~x[17] & ~x[18];
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & x[48];
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & x[10] & x[13];
			partial_clause[5][91] 	= partial_clause_prev[5][91] & x[33];
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & x[21];
			partial_clause[5][95] 	= partial_clause_prev[5][95] & ~x[42] & ~x[44];
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & ~x[12] & ~x[13] & ~x[44];
			partial_clause[5][99] 	= partial_clause_prev[5][99] & x[21];
			partial_clause[5][100] 	= partial_clause_prev[5][100] & 1'b1;
			partial_clause[5][101] 	= partial_clause_prev[5][101] & 1'b1;
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & x[46];
			partial_clause[5][104] 	= partial_clause_prev[5][104] & 1'b1;
			partial_clause[5][105] 	= partial_clause_prev[5][105] & 1'b1;
			partial_clause[5][106] 	= partial_clause_prev[5][106] & x[23];
			partial_clause[5][107] 	= partial_clause_prev[5][107] & 1'b1;
			partial_clause[5][108] 	= partial_clause_prev[5][108] & 1'b1;
			partial_clause[5][109] 	= partial_clause_prev[5][109] & x[13] & ~x[17] & x[41] & ~x[44];
			partial_clause[5][110] 	= partial_clause_prev[5][110] & ~x[10] & x[13];
			partial_clause[5][111] 	= partial_clause_prev[5][111] & 1'b1;
			partial_clause[5][112] 	= partial_clause_prev[5][112] & x[26];
			partial_clause[5][113] 	= partial_clause_prev[5][113] & 1'b1;
			partial_clause[5][114] 	= partial_clause_prev[5][114] & 1'b1;
			partial_clause[5][115] 	= partial_clause_prev[5][115] & 1'b1;
			partial_clause[5][116] 	= partial_clause_prev[5][116] & 1'b1;
			partial_clause[5][117] 	= partial_clause_prev[5][117] & 1'b1;
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & x[0];
			partial_clause[5][120] 	= partial_clause_prev[5][120] & 1'b1;
			partial_clause[5][121] 	= partial_clause_prev[5][121] & x[44];
			partial_clause[5][122] 	= partial_clause_prev[5][122] & ~x[13];
			partial_clause[5][123] 	= partial_clause_prev[5][123] & x[28];
			partial_clause[5][124] 	= partial_clause_prev[5][124] & 1'b1;
			partial_clause[5][125] 	= partial_clause_prev[5][125] & 1'b1;
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & 1'b1;
			partial_clause[5][128] 	= partial_clause_prev[5][128] & 1'b1;
			partial_clause[5][129] 	= partial_clause_prev[5][129] & 1'b1;
			partial_clause[5][130] 	= partial_clause_prev[5][130] & 1'b1;
			partial_clause[5][131] 	= partial_clause_prev[5][131] & 1'b1;
			partial_clause[5][132] 	= partial_clause_prev[5][132] & ~x[17];
			partial_clause[5][133] 	= partial_clause_prev[5][133] & x[27];
			partial_clause[5][134] 	= partial_clause_prev[5][134] & 1'b1;
			partial_clause[5][135] 	= partial_clause_prev[5][135] & 1'b1;
			partial_clause[5][136] 	= partial_clause_prev[5][136] & x[16];
			partial_clause[5][137] 	= partial_clause_prev[5][137] & 1'b1;
			partial_clause[5][138] 	= partial_clause_prev[5][138] & 1'b1;
			partial_clause[5][139] 	= partial_clause_prev[5][139] & 1'b1;
			partial_clause[5][140] 	= partial_clause_prev[5][140] & 1'b1;
			partial_clause[5][141] 	= partial_clause_prev[5][141] & 1'b1;
			partial_clause[5][142] 	= partial_clause_prev[5][142] & 1'b1;
			partial_clause[5][143] 	= partial_clause_prev[5][143] & x[14] & ~x[38];
			partial_clause[5][144] 	= partial_clause_prev[5][144] & 1'b1;
			partial_clause[5][145] 	= partial_clause_prev[5][145] & 1'b1;
			partial_clause[5][146] 	= partial_clause_prev[5][146] & 1'b1;
			partial_clause[5][147] 	= partial_clause_prev[5][147] & x[13];
			partial_clause[5][148] 	= partial_clause_prev[5][148] & x[43];
			partial_clause[5][149] 	= partial_clause_prev[5][149] & x[0];
			partial_clause[5][150] 	= partial_clause_prev[5][150] & 1'b1;
			partial_clause[5][151] 	= partial_clause_prev[5][151] & 1'b1;
			partial_clause[5][152] 	= partial_clause_prev[5][152] & ~x[19] & ~x[35];
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & 1'b1;
			partial_clause[5][155] 	= partial_clause_prev[5][155] & 1'b1;
			partial_clause[5][156] 	= partial_clause_prev[5][156] & x[44];
			partial_clause[5][157] 	= partial_clause_prev[5][157] & 1'b1;
			partial_clause[5][158] 	= partial_clause_prev[5][158] & 1'b1;
			partial_clause[5][159] 	= partial_clause_prev[5][159] & 1'b1;
			partial_clause[5][160] 	= partial_clause_prev[5][160] & 1'b1;
			partial_clause[5][161] 	= partial_clause_prev[5][161] & 1'b1;
			partial_clause[5][162] 	= partial_clause_prev[5][162] & 1'b1;
			partial_clause[5][163] 	= partial_clause_prev[5][163] & 1'b1;
			partial_clause[5][164] 	= partial_clause_prev[5][164] & ~x[63];
			partial_clause[5][165] 	= partial_clause_prev[5][165] & 1'b1;
			partial_clause[5][166] 	= partial_clause_prev[5][166] & 1'b1;
			partial_clause[5][167] 	= partial_clause_prev[5][167] & 1'b1;
			partial_clause[5][168] 	= partial_clause_prev[5][168] & 1'b1;
			partial_clause[5][169] 	= partial_clause_prev[5][169] & ~x[48];
			partial_clause[5][170] 	= partial_clause_prev[5][170] & 1'b1;
			partial_clause[5][171] 	= partial_clause_prev[5][171] & 1'b1;
			partial_clause[5][172] 	= partial_clause_prev[5][172] & 1'b1;
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & 1'b1;
			partial_clause[5][175] 	= partial_clause_prev[5][175] & 1'b1;
			partial_clause[5][176] 	= partial_clause_prev[5][176] & 1'b1;
			partial_clause[5][177] 	= partial_clause_prev[5][177] & ~x[49];
			partial_clause[5][178] 	= partial_clause_prev[5][178] & 1'b1;
			partial_clause[5][179] 	= partial_clause_prev[5][179] & ~x[63];
			partial_clause[5][180] 	= partial_clause_prev[5][180] & 1'b1;
			partial_clause[5][181] 	= partial_clause_prev[5][181] & ~x[7] & ~x[17] & ~x[59] & ~x[61];
			partial_clause[5][182] 	= partial_clause_prev[5][182] & 1'b1;
			partial_clause[5][183] 	= partial_clause_prev[5][183] & 1'b1;
			partial_clause[5][184] 	= partial_clause_prev[5][184] & 1'b1;
			partial_clause[5][185] 	= partial_clause_prev[5][185] & 1'b1;
			partial_clause[5][186] 	= partial_clause_prev[5][186] & x[41] & ~x[45];
			partial_clause[5][187] 	= partial_clause_prev[5][187] & 1'b1;
			partial_clause[5][188] 	= partial_clause_prev[5][188] & 1'b1;
			partial_clause[5][189] 	= partial_clause_prev[5][189] & ~x[19] & x[40] & ~x[48];
			partial_clause[5][190] 	= partial_clause_prev[5][190] & 1'b1;
			partial_clause[5][191] 	= partial_clause_prev[5][191] & 1'b1;
			partial_clause[5][192] 	= partial_clause_prev[5][192] & 1'b1;
			partial_clause[5][193] 	= partial_clause_prev[5][193] & ~x[47];
			partial_clause[5][194] 	= partial_clause_prev[5][194] & 1'b1;
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & 1'b1;
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & 1'b1;
			partial_clause[5][199] 	= partial_clause_prev[5][199] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & ~x[43] & x[62];
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & ~x[41];
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & ~x[17] & ~x[42];
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & ~x[11] & ~x[38];
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & ~x[9];
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & ~x[44];
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & ~x[14];
			partial_clause[6][22] 	= partial_clause_prev[6][22] & ~x[8] & ~x[55];
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & ~x[14] & ~x[18] & ~x[41];
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & ~x[10];
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & ~x[61];
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & ~x[7];
			partial_clause[6][42] 	= partial_clause_prev[6][42] & ~x[11] & ~x[38];
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & ~x[17];
			partial_clause[6][46] 	= partial_clause_prev[6][46] & ~x[45];
			partial_clause[6][47] 	= partial_clause_prev[6][47] & x[11];
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & ~x[13] & ~x[15];
			partial_clause[6][53] 	= partial_clause_prev[6][53] & ~x[16] & ~x[19] & ~x[41] & ~x[45];
			partial_clause[6][54] 	= partial_clause_prev[6][54] & ~x[14] & x[36];
			partial_clause[6][55] 	= partial_clause_prev[6][55] & x[9];
			partial_clause[6][56] 	= partial_clause_prev[6][56] & ~x[39];
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & ~x[46];
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & ~x[46];
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & ~x[10] & ~x[12];
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & ~x[63];
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & ~x[9];
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & ~x[12];
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & ~x[12];
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & ~x[9] & ~x[37];
			partial_clause[6][94] 	= partial_clause_prev[6][94] & x[12];
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			partial_clause[6][100] 	= partial_clause_prev[6][100] & 1'b1;
			partial_clause[6][101] 	= partial_clause_prev[6][101] & x[17];
			partial_clause[6][102] 	= partial_clause_prev[6][102] & x[42];
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & 1'b1;
			partial_clause[6][105] 	= partial_clause_prev[6][105] & 1'b1;
			partial_clause[6][106] 	= partial_clause_prev[6][106] & ~x[45];
			partial_clause[6][107] 	= partial_clause_prev[6][107] & x[41];
			partial_clause[6][108] 	= partial_clause_prev[6][108] & 1'b1;
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & x[15];
			partial_clause[6][111] 	= partial_clause_prev[6][111] & 1'b1;
			partial_clause[6][112] 	= partial_clause_prev[6][112] & 1'b1;
			partial_clause[6][113] 	= partial_clause_prev[6][113] & x[15];
			partial_clause[6][114] 	= partial_clause_prev[6][114] & 1'b1;
			partial_clause[6][115] 	= partial_clause_prev[6][115] & x[39];
			partial_clause[6][116] 	= partial_clause_prev[6][116] & 1'b1;
			partial_clause[6][117] 	= partial_clause_prev[6][117] & 1'b1;
			partial_clause[6][118] 	= partial_clause_prev[6][118] & x[12];
			partial_clause[6][119] 	= partial_clause_prev[6][119] & 1'b1;
			partial_clause[6][120] 	= partial_clause_prev[6][120] & 1'b1;
			partial_clause[6][121] 	= partial_clause_prev[6][121] & 1'b1;
			partial_clause[6][122] 	= partial_clause_prev[6][122] & x[41];
			partial_clause[6][123] 	= partial_clause_prev[6][123] & 1'b1;
			partial_clause[6][124] 	= partial_clause_prev[6][124] & 1'b1;
			partial_clause[6][125] 	= partial_clause_prev[6][125] & ~x[46];
			partial_clause[6][126] 	= partial_clause_prev[6][126] & x[13];
			partial_clause[6][127] 	= partial_clause_prev[6][127] & 1'b1;
			partial_clause[6][128] 	= partial_clause_prev[6][128] & 1'b1;
			partial_clause[6][129] 	= partial_clause_prev[6][129] & 1'b1;
			partial_clause[6][130] 	= partial_clause_prev[6][130] & x[16];
			partial_clause[6][131] 	= partial_clause_prev[6][131] & 1'b1;
			partial_clause[6][132] 	= partial_clause_prev[6][132] & x[20];
			partial_clause[6][133] 	= partial_clause_prev[6][133] & 1'b1;
			partial_clause[6][134] 	= partial_clause_prev[6][134] & x[43];
			partial_clause[6][135] 	= partial_clause_prev[6][135] & 1'b1;
			partial_clause[6][136] 	= partial_clause_prev[6][136] & ~x[39];
			partial_clause[6][137] 	= partial_clause_prev[6][137] & x[43];
			partial_clause[6][138] 	= partial_clause_prev[6][138] & x[18];
			partial_clause[6][139] 	= partial_clause_prev[6][139] & x[12];
			partial_clause[6][140] 	= partial_clause_prev[6][140] & x[42];
			partial_clause[6][141] 	= partial_clause_prev[6][141] & 1'b1;
			partial_clause[6][142] 	= partial_clause_prev[6][142] & 1'b1;
			partial_clause[6][143] 	= partial_clause_prev[6][143] & x[40];
			partial_clause[6][144] 	= partial_clause_prev[6][144] & 1'b1;
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & 1'b1;
			partial_clause[6][147] 	= partial_clause_prev[6][147] & x[19];
			partial_clause[6][148] 	= partial_clause_prev[6][148] & 1'b1;
			partial_clause[6][149] 	= partial_clause_prev[6][149] & 1'b1;
			partial_clause[6][150] 	= partial_clause_prev[6][150] & 1'b1;
			partial_clause[6][151] 	= partial_clause_prev[6][151] & 1'b1;
			partial_clause[6][152] 	= partial_clause_prev[6][152] & 1'b1;
			partial_clause[6][153] 	= partial_clause_prev[6][153] & 1'b1;
			partial_clause[6][154] 	= partial_clause_prev[6][154] & 1'b1;
			partial_clause[6][155] 	= partial_clause_prev[6][155] & 1'b1;
			partial_clause[6][156] 	= partial_clause_prev[6][156] & x[13];
			partial_clause[6][157] 	= partial_clause_prev[6][157] & 1'b1;
			partial_clause[6][158] 	= partial_clause_prev[6][158] & 1'b1;
			partial_clause[6][159] 	= partial_clause_prev[6][159] & 1'b1;
			partial_clause[6][160] 	= partial_clause_prev[6][160] & 1'b1;
			partial_clause[6][161] 	= partial_clause_prev[6][161] & 1'b1;
			partial_clause[6][162] 	= partial_clause_prev[6][162] & 1'b1;
			partial_clause[6][163] 	= partial_clause_prev[6][163] & 1'b1;
			partial_clause[6][164] 	= partial_clause_prev[6][164] & 1'b1;
			partial_clause[6][165] 	= partial_clause_prev[6][165] & x[19];
			partial_clause[6][166] 	= partial_clause_prev[6][166] & x[16];
			partial_clause[6][167] 	= partial_clause_prev[6][167] & 1'b1;
			partial_clause[6][168] 	= partial_clause_prev[6][168] & 1'b1;
			partial_clause[6][169] 	= partial_clause_prev[6][169] & 1'b1;
			partial_clause[6][170] 	= partial_clause_prev[6][170] & 1'b1;
			partial_clause[6][171] 	= partial_clause_prev[6][171] & 1'b1;
			partial_clause[6][172] 	= partial_clause_prev[6][172] & 1'b1;
			partial_clause[6][173] 	= partial_clause_prev[6][173] & 1'b1;
			partial_clause[6][174] 	= partial_clause_prev[6][174] & 1'b1;
			partial_clause[6][175] 	= partial_clause_prev[6][175] & 1'b1;
			partial_clause[6][176] 	= partial_clause_prev[6][176] & ~x[33] & ~x[34];
			partial_clause[6][177] 	= partial_clause_prev[6][177] & 1'b1;
			partial_clause[6][178] 	= partial_clause_prev[6][178] & 1'b1;
			partial_clause[6][179] 	= partial_clause_prev[6][179] & x[45];
			partial_clause[6][180] 	= partial_clause_prev[6][180] & 1'b1;
			partial_clause[6][181] 	= partial_clause_prev[6][181] & 1'b1;
			partial_clause[6][182] 	= partial_clause_prev[6][182] & 1'b1;
			partial_clause[6][183] 	= partial_clause_prev[6][183] & 1'b1;
			partial_clause[6][184] 	= partial_clause_prev[6][184] & 1'b1;
			partial_clause[6][185] 	= partial_clause_prev[6][185] & 1'b1;
			partial_clause[6][186] 	= partial_clause_prev[6][186] & x[39];
			partial_clause[6][187] 	= partial_clause_prev[6][187] & x[14];
			partial_clause[6][188] 	= partial_clause_prev[6][188] & 1'b1;
			partial_clause[6][189] 	= partial_clause_prev[6][189] & 1'b1;
			partial_clause[6][190] 	= partial_clause_prev[6][190] & 1'b1;
			partial_clause[6][191] 	= partial_clause_prev[6][191] & 1'b1;
			partial_clause[6][192] 	= partial_clause_prev[6][192] & 1'b1;
			partial_clause[6][193] 	= partial_clause_prev[6][193] & 1'b1;
			partial_clause[6][194] 	= partial_clause_prev[6][194] & 1'b1;
			partial_clause[6][195] 	= partial_clause_prev[6][195] & 1'b1;
			partial_clause[6][196] 	= partial_clause_prev[6][196] & 1'b1;
			partial_clause[6][197] 	= partial_clause_prev[6][197] & 1'b1;
			partial_clause[6][198] 	= partial_clause_prev[6][198] & 1'b1;
			partial_clause[6][199] 	= partial_clause_prev[6][199] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & x[8] & x[39];
			partial_clause[7][1] 	= partial_clause_prev[7][1] & x[42];
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & x[54];
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & x[1];
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & x[7];
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & x[55];
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & x[37] & x[39];
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & x[1];
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & x[12];
			partial_clause[7][42] 	= partial_clause_prev[7][42] & x[41];
			partial_clause[7][43] 	= partial_clause_prev[7][43] & x[0];
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & x[10] & x[40];
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & ~x[60] & ~x[63];
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & x[35] & x[37];
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & ~x[30];
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & x[4] & x[8];
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & x[29];
			partial_clause[7][100] 	= partial_clause_prev[7][100] & 1'b1;
			partial_clause[7][101] 	= partial_clause_prev[7][101] & 1'b1;
			partial_clause[7][102] 	= partial_clause_prev[7][102] & 1'b1;
			partial_clause[7][103] 	= partial_clause_prev[7][103] & 1'b1;
			partial_clause[7][104] 	= partial_clause_prev[7][104] & ~x[2];
			partial_clause[7][105] 	= partial_clause_prev[7][105] & ~x[10];
			partial_clause[7][106] 	= partial_clause_prev[7][106] & 1'b1;
			partial_clause[7][107] 	= partial_clause_prev[7][107] & 1'b1;
			partial_clause[7][108] 	= partial_clause_prev[7][108] & ~x[8];
			partial_clause[7][109] 	= partial_clause_prev[7][109] & ~x[5] & ~x[61];
			partial_clause[7][110] 	= partial_clause_prev[7][110] & 1'b1;
			partial_clause[7][111] 	= partial_clause_prev[7][111] & 1'b1;
			partial_clause[7][112] 	= partial_clause_prev[7][112] & 1'b1;
			partial_clause[7][113] 	= partial_clause_prev[7][113] & ~x[61];
			partial_clause[7][114] 	= partial_clause_prev[7][114] & 1'b1;
			partial_clause[7][115] 	= partial_clause_prev[7][115] & 1'b1;
			partial_clause[7][116] 	= partial_clause_prev[7][116] & 1'b1;
			partial_clause[7][117] 	= partial_clause_prev[7][117] & 1'b1;
			partial_clause[7][118] 	= partial_clause_prev[7][118] & 1'b1;
			partial_clause[7][119] 	= partial_clause_prev[7][119] & 1'b1;
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & 1'b1;
			partial_clause[7][123] 	= partial_clause_prev[7][123] & 1'b1;
			partial_clause[7][124] 	= partial_clause_prev[7][124] & 1'b1;
			partial_clause[7][125] 	= partial_clause_prev[7][125] & 1'b1;
			partial_clause[7][126] 	= partial_clause_prev[7][126] & 1'b1;
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & 1'b1;
			partial_clause[7][129] 	= partial_clause_prev[7][129] & 1'b1;
			partial_clause[7][130] 	= partial_clause_prev[7][130] & ~x[2] & ~x[12];
			partial_clause[7][131] 	= partial_clause_prev[7][131] & 1'b1;
			partial_clause[7][132] 	= partial_clause_prev[7][132] & 1'b1;
			partial_clause[7][133] 	= partial_clause_prev[7][133] & 1'b1;
			partial_clause[7][134] 	= partial_clause_prev[7][134] & 1'b1;
			partial_clause[7][135] 	= partial_clause_prev[7][135] & 1'b1;
			partial_clause[7][136] 	= partial_clause_prev[7][136] & ~x[40];
			partial_clause[7][137] 	= partial_clause_prev[7][137] & ~x[30] & ~x[43];
			partial_clause[7][138] 	= partial_clause_prev[7][138] & 1'b1;
			partial_clause[7][139] 	= partial_clause_prev[7][139] & 1'b1;
			partial_clause[7][140] 	= partial_clause_prev[7][140] & 1'b1;
			partial_clause[7][141] 	= partial_clause_prev[7][141] & ~x[5] & ~x[60];
			partial_clause[7][142] 	= partial_clause_prev[7][142] & 1'b1;
			partial_clause[7][143] 	= partial_clause_prev[7][143] & 1'b1;
			partial_clause[7][144] 	= partial_clause_prev[7][144] & 1'b1;
			partial_clause[7][145] 	= partial_clause_prev[7][145] & 1'b1;
			partial_clause[7][146] 	= partial_clause_prev[7][146] & 1'b1;
			partial_clause[7][147] 	= partial_clause_prev[7][147] & 1'b1;
			partial_clause[7][148] 	= partial_clause_prev[7][148] & 1'b1;
			partial_clause[7][149] 	= partial_clause_prev[7][149] & 1'b1;
			partial_clause[7][150] 	= partial_clause_prev[7][150] & 1'b1;
			partial_clause[7][151] 	= partial_clause_prev[7][151] & 1'b1;
			partial_clause[7][152] 	= partial_clause_prev[7][152] & 1'b1;
			partial_clause[7][153] 	= partial_clause_prev[7][153] & 1'b1;
			partial_clause[7][154] 	= partial_clause_prev[7][154] & 1'b1;
			partial_clause[7][155] 	= partial_clause_prev[7][155] & 1'b1;
			partial_clause[7][156] 	= partial_clause_prev[7][156] & 1'b1;
			partial_clause[7][157] 	= partial_clause_prev[7][157] & ~x[11];
			partial_clause[7][158] 	= partial_clause_prev[7][158] & 1'b1;
			partial_clause[7][159] 	= partial_clause_prev[7][159] & ~x[13] & ~x[41];
			partial_clause[7][160] 	= partial_clause_prev[7][160] & 1'b1;
			partial_clause[7][161] 	= partial_clause_prev[7][161] & 1'b1;
			partial_clause[7][162] 	= partial_clause_prev[7][162] & 1'b1;
			partial_clause[7][163] 	= partial_clause_prev[7][163] & ~x[39];
			partial_clause[7][164] 	= partial_clause_prev[7][164] & 1'b1;
			partial_clause[7][165] 	= partial_clause_prev[7][165] & 1'b1;
			partial_clause[7][166] 	= partial_clause_prev[7][166] & 1'b1;
			partial_clause[7][167] 	= partial_clause_prev[7][167] & 1'b1;
			partial_clause[7][168] 	= partial_clause_prev[7][168] & 1'b1;
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & 1'b1;
			partial_clause[7][171] 	= partial_clause_prev[7][171] & 1'b1;
			partial_clause[7][172] 	= partial_clause_prev[7][172] & 1'b1;
			partial_clause[7][173] 	= partial_clause_prev[7][173] & 1'b1;
			partial_clause[7][174] 	= partial_clause_prev[7][174] & 1'b1;
			partial_clause[7][175] 	= partial_clause_prev[7][175] & 1'b1;
			partial_clause[7][176] 	= partial_clause_prev[7][176] & 1'b1;
			partial_clause[7][177] 	= partial_clause_prev[7][177] & 1'b1;
			partial_clause[7][178] 	= partial_clause_prev[7][178] & 1'b1;
			partial_clause[7][179] 	= partial_clause_prev[7][179] & 1'b1;
			partial_clause[7][180] 	= partial_clause_prev[7][180] & 1'b1;
			partial_clause[7][181] 	= partial_clause_prev[7][181] & 1'b1;
			partial_clause[7][182] 	= partial_clause_prev[7][182] & 1'b1;
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & 1'b1;
			partial_clause[7][185] 	= partial_clause_prev[7][185] & 1'b1;
			partial_clause[7][186] 	= partial_clause_prev[7][186] & ~x[43];
			partial_clause[7][187] 	= partial_clause_prev[7][187] & 1'b1;
			partial_clause[7][188] 	= partial_clause_prev[7][188] & 1'b1;
			partial_clause[7][189] 	= partial_clause_prev[7][189] & 1'b1;
			partial_clause[7][190] 	= partial_clause_prev[7][190] & 1'b1;
			partial_clause[7][191] 	= partial_clause_prev[7][191] & 1'b1;
			partial_clause[7][192] 	= partial_clause_prev[7][192] & 1'b1;
			partial_clause[7][193] 	= partial_clause_prev[7][193] & ~x[5] & ~x[14];
			partial_clause[7][194] 	= partial_clause_prev[7][194] & 1'b1;
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & 1'b1;
			partial_clause[7][197] 	= partial_clause_prev[7][197] & 1'b1;
			partial_clause[7][198] 	= partial_clause_prev[7][198] & ~x[60];
			partial_clause[7][199] 	= partial_clause_prev[7][199] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & ~x[40];
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & x[18];
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & x[62];
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & ~x[40];
			partial_clause[8][19] 	= partial_clause_prev[8][19] & ~x[42];
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & ~x[11];
			partial_clause[8][22] 	= partial_clause_prev[8][22] & ~x[11];
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & x[58];
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & ~x[11];
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & x[57];
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & x[44];
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & ~x[40];
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & x[63];
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & ~x[40];
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & x[63];
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & x[47];
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & x[33];
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & x[22];
			partial_clause[8][73] 	= partial_clause_prev[8][73] & x[47];
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & x[57];
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & x[61];
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & x[31];
			partial_clause[8][84] 	= partial_clause_prev[8][84] & x[50];
			partial_clause[8][85] 	= partial_clause_prev[8][85] & x[37];
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & x[32] & ~x[35];
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			partial_clause[8][100] 	= partial_clause_prev[8][100] & 1'b1;
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & 1'b1;
			partial_clause[8][103] 	= partial_clause_prev[8][103] & 1'b1;
			partial_clause[8][104] 	= partial_clause_prev[8][104] & 1'b1;
			partial_clause[8][105] 	= partial_clause_prev[8][105] & 1'b1;
			partial_clause[8][106] 	= partial_clause_prev[8][106] & 1'b1;
			partial_clause[8][107] 	= partial_clause_prev[8][107] & 1'b1;
			partial_clause[8][108] 	= partial_clause_prev[8][108] & 1'b1;
			partial_clause[8][109] 	= partial_clause_prev[8][109] & 1'b1;
			partial_clause[8][110] 	= partial_clause_prev[8][110] & 1'b1;
			partial_clause[8][111] 	= partial_clause_prev[8][111] & 1'b1;
			partial_clause[8][112] 	= partial_clause_prev[8][112] & 1'b1;
			partial_clause[8][113] 	= partial_clause_prev[8][113] & ~x[46];
			partial_clause[8][114] 	= partial_clause_prev[8][114] & 1'b1;
			partial_clause[8][115] 	= partial_clause_prev[8][115] & 1'b1;
			partial_clause[8][116] 	= partial_clause_prev[8][116] & 1'b1;
			partial_clause[8][117] 	= partial_clause_prev[8][117] & 1'b1;
			partial_clause[8][118] 	= partial_clause_prev[8][118] & 1'b1;
			partial_clause[8][119] 	= partial_clause_prev[8][119] & 1'b1;
			partial_clause[8][120] 	= partial_clause_prev[8][120] & 1'b1;
			partial_clause[8][121] 	= partial_clause_prev[8][121] & 1'b1;
			partial_clause[8][122] 	= partial_clause_prev[8][122] & 1'b1;
			partial_clause[8][123] 	= partial_clause_prev[8][123] & 1'b1;
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & 1'b1;
			partial_clause[8][126] 	= partial_clause_prev[8][126] & 1'b1;
			partial_clause[8][127] 	= partial_clause_prev[8][127] & ~x[21];
			partial_clause[8][128] 	= partial_clause_prev[8][128] & 1'b1;
			partial_clause[8][129] 	= partial_clause_prev[8][129] & 1'b1;
			partial_clause[8][130] 	= partial_clause_prev[8][130] & 1'b1;
			partial_clause[8][131] 	= partial_clause_prev[8][131] & 1'b1;
			partial_clause[8][132] 	= partial_clause_prev[8][132] & 1'b1;
			partial_clause[8][133] 	= partial_clause_prev[8][133] & ~x[9] & ~x[36] & ~x[47] & ~x[62];
			partial_clause[8][134] 	= partial_clause_prev[8][134] & 1'b1;
			partial_clause[8][135] 	= partial_clause_prev[8][135] & 1'b1;
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & 1'b1;
			partial_clause[8][138] 	= partial_clause_prev[8][138] & 1'b1;
			partial_clause[8][139] 	= partial_clause_prev[8][139] & 1'b1;
			partial_clause[8][140] 	= partial_clause_prev[8][140] & 1'b1;
			partial_clause[8][141] 	= partial_clause_prev[8][141] & ~x[18];
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & 1'b1;
			partial_clause[8][144] 	= partial_clause_prev[8][144] & 1'b1;
			partial_clause[8][145] 	= partial_clause_prev[8][145] & ~x[6] & ~x[8] & ~x[15];
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & 1'b1;
			partial_clause[8][148] 	= partial_clause_prev[8][148] & 1'b1;
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & 1'b1;
			partial_clause[8][151] 	= partial_clause_prev[8][151] & 1'b1;
			partial_clause[8][152] 	= partial_clause_prev[8][152] & 1'b1;
			partial_clause[8][153] 	= partial_clause_prev[8][153] & ~x[47];
			partial_clause[8][154] 	= partial_clause_prev[8][154] & 1'b1;
			partial_clause[8][155] 	= partial_clause_prev[8][155] & 1'b1;
			partial_clause[8][156] 	= partial_clause_prev[8][156] & 1'b1;
			partial_clause[8][157] 	= partial_clause_prev[8][157] & 1'b1;
			partial_clause[8][158] 	= partial_clause_prev[8][158] & 1'b1;
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & 1'b1;
			partial_clause[8][161] 	= partial_clause_prev[8][161] & 1'b1;
			partial_clause[8][162] 	= partial_clause_prev[8][162] & 1'b1;
			partial_clause[8][163] 	= partial_clause_prev[8][163] & 1'b1;
			partial_clause[8][164] 	= partial_clause_prev[8][164] & ~x[36];
			partial_clause[8][165] 	= partial_clause_prev[8][165] & ~x[47];
			partial_clause[8][166] 	= partial_clause_prev[8][166] & 1'b1;
			partial_clause[8][167] 	= partial_clause_prev[8][167] & 1'b1;
			partial_clause[8][168] 	= partial_clause_prev[8][168] & 1'b1;
			partial_clause[8][169] 	= partial_clause_prev[8][169] & ~x[9] & ~x[33] & ~x[34] & ~x[35] & ~x[60];
			partial_clause[8][170] 	= partial_clause_prev[8][170] & 1'b1;
			partial_clause[8][171] 	= partial_clause_prev[8][171] & 1'b1;
			partial_clause[8][172] 	= partial_clause_prev[8][172] & 1'b1;
			partial_clause[8][173] 	= partial_clause_prev[8][173] & 1'b1;
			partial_clause[8][174] 	= partial_clause_prev[8][174] & 1'b1;
			partial_clause[8][175] 	= partial_clause_prev[8][175] & 1'b1;
			partial_clause[8][176] 	= partial_clause_prev[8][176] & 1'b1;
			partial_clause[8][177] 	= partial_clause_prev[8][177] & 1'b1;
			partial_clause[8][178] 	= partial_clause_prev[8][178] & 1'b1;
			partial_clause[8][179] 	= partial_clause_prev[8][179] & 1'b1;
			partial_clause[8][180] 	= partial_clause_prev[8][180] & 1'b1;
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & ~x[8] & ~x[61];
			partial_clause[8][183] 	= partial_clause_prev[8][183] & ~x[20];
			partial_clause[8][184] 	= partial_clause_prev[8][184] & 1'b1;
			partial_clause[8][185] 	= partial_clause_prev[8][185] & 1'b1;
			partial_clause[8][186] 	= partial_clause_prev[8][186] & 1'b1;
			partial_clause[8][187] 	= partial_clause_prev[8][187] & 1'b1;
			partial_clause[8][188] 	= partial_clause_prev[8][188] & 1'b1;
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & 1'b1;
			partial_clause[8][191] 	= partial_clause_prev[8][191] & 1'b1;
			partial_clause[8][192] 	= partial_clause_prev[8][192] & 1'b1;
			partial_clause[8][193] 	= partial_clause_prev[8][193] & 1'b1;
			partial_clause[8][194] 	= partial_clause_prev[8][194] & 1'b1;
			partial_clause[8][195] 	= partial_clause_prev[8][195] & 1'b1;
			partial_clause[8][196] 	= partial_clause_prev[8][196] & 1'b1;
			partial_clause[8][197] 	= partial_clause_prev[8][197] & 1'b1;
			partial_clause[8][198] 	= partial_clause_prev[8][198] & 1'b1;
			partial_clause[8][199] 	= partial_clause_prev[8][199] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & ~x[37];
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & x[61];
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & ~x[36];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & ~x[5] & x[35];
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & ~x[3];
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & ~x[4];
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & ~x[4] & x[8];
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & ~x[2] & ~x[3];
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & ~x[37] & ~x[38];
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
			partial_clause[9][100] 	= partial_clause_prev[9][100] & 1'b1;
			partial_clause[9][101] 	= partial_clause_prev[9][101] & 1'b1;
			partial_clause[9][102] 	= partial_clause_prev[9][102] & 1'b1;
			partial_clause[9][103] 	= partial_clause_prev[9][103] & 1'b1;
			partial_clause[9][104] 	= partial_clause_prev[9][104] & 1'b1;
			partial_clause[9][105] 	= partial_clause_prev[9][105] & 1'b1;
			partial_clause[9][106] 	= partial_clause_prev[9][106] & 1'b1;
			partial_clause[9][107] 	= partial_clause_prev[9][107] & 1'b1;
			partial_clause[9][108] 	= partial_clause_prev[9][108] & 1'b1;
			partial_clause[9][109] 	= partial_clause_prev[9][109] & ~x[10];
			partial_clause[9][110] 	= partial_clause_prev[9][110] & 1'b1;
			partial_clause[9][111] 	= partial_clause_prev[9][111] & ~x[63];
			partial_clause[9][112] 	= partial_clause_prev[9][112] & 1'b1;
			partial_clause[9][113] 	= partial_clause_prev[9][113] & ~x[11] & ~x[12];
			partial_clause[9][114] 	= partial_clause_prev[9][114] & 1'b1;
			partial_clause[9][115] 	= partial_clause_prev[9][115] & 1'b1;
			partial_clause[9][116] 	= partial_clause_prev[9][116] & 1'b1;
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & 1'b1;
			partial_clause[9][119] 	= partial_clause_prev[9][119] & ~x[35] & ~x[36] & ~x[61];
			partial_clause[9][120] 	= partial_clause_prev[9][120] & 1'b1;
			partial_clause[9][121] 	= partial_clause_prev[9][121] & 1'b1;
			partial_clause[9][122] 	= partial_clause_prev[9][122] & 1'b1;
			partial_clause[9][123] 	= partial_clause_prev[9][123] & 1'b1;
			partial_clause[9][124] 	= partial_clause_prev[9][124] & ~x[59];
			partial_clause[9][125] 	= partial_clause_prev[9][125] & 1'b1;
			partial_clause[9][126] 	= partial_clause_prev[9][126] & 1'b1;
			partial_clause[9][127] 	= partial_clause_prev[9][127] & 1'b1;
			partial_clause[9][128] 	= partial_clause_prev[9][128] & 1'b1;
			partial_clause[9][129] 	= partial_clause_prev[9][129] & 1'b1;
			partial_clause[9][130] 	= partial_clause_prev[9][130] & 1'b1;
			partial_clause[9][131] 	= partial_clause_prev[9][131] & 1'b1;
			partial_clause[9][132] 	= partial_clause_prev[9][132] & 1'b1;
			partial_clause[9][133] 	= partial_clause_prev[9][133] & 1'b1;
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & 1'b1;
			partial_clause[9][138] 	= partial_clause_prev[9][138] & 1'b1;
			partial_clause[9][139] 	= partial_clause_prev[9][139] & 1'b1;
			partial_clause[9][140] 	= partial_clause_prev[9][140] & 1'b1;
			partial_clause[9][141] 	= partial_clause_prev[9][141] & 1'b1;
			partial_clause[9][142] 	= partial_clause_prev[9][142] & 1'b1;
			partial_clause[9][143] 	= partial_clause_prev[9][143] & 1'b1;
			partial_clause[9][144] 	= partial_clause_prev[9][144] & 1'b1;
			partial_clause[9][145] 	= partial_clause_prev[9][145] & 1'b1;
			partial_clause[9][146] 	= partial_clause_prev[9][146] & 1'b1;
			partial_clause[9][147] 	= partial_clause_prev[9][147] & ~x[61] & ~x[63];
			partial_clause[9][148] 	= partial_clause_prev[9][148] & 1'b1;
			partial_clause[9][149] 	= partial_clause_prev[9][149] & 1'b1;
			partial_clause[9][150] 	= partial_clause_prev[9][150] & 1'b1;
			partial_clause[9][151] 	= partial_clause_prev[9][151] & 1'b1;
			partial_clause[9][152] 	= partial_clause_prev[9][152] & 1'b1;
			partial_clause[9][153] 	= partial_clause_prev[9][153] & 1'b1;
			partial_clause[9][154] 	= partial_clause_prev[9][154] & 1'b1;
			partial_clause[9][155] 	= partial_clause_prev[9][155] & 1'b1;
			partial_clause[9][156] 	= partial_clause_prev[9][156] & 1'b1;
			partial_clause[9][157] 	= partial_clause_prev[9][157] & 1'b1;
			partial_clause[9][158] 	= partial_clause_prev[9][158] & 1'b1;
			partial_clause[9][159] 	= partial_clause_prev[9][159] & 1'b1;
			partial_clause[9][160] 	= partial_clause_prev[9][160] & 1'b1;
			partial_clause[9][161] 	= partial_clause_prev[9][161] & 1'b1;
			partial_clause[9][162] 	= partial_clause_prev[9][162] & 1'b1;
			partial_clause[9][163] 	= partial_clause_prev[9][163] & 1'b1;
			partial_clause[9][164] 	= partial_clause_prev[9][164] & 1'b1;
			partial_clause[9][165] 	= partial_clause_prev[9][165] & 1'b1;
			partial_clause[9][166] 	= partial_clause_prev[9][166] & 1'b1;
			partial_clause[9][167] 	= partial_clause_prev[9][167] & 1'b1;
			partial_clause[9][168] 	= partial_clause_prev[9][168] & 1'b1;
			partial_clause[9][169] 	= partial_clause_prev[9][169] & 1'b1;
			partial_clause[9][170] 	= partial_clause_prev[9][170] & 1'b1;
			partial_clause[9][171] 	= partial_clause_prev[9][171] & 1'b1;
			partial_clause[9][172] 	= partial_clause_prev[9][172] & 1'b1;
			partial_clause[9][173] 	= partial_clause_prev[9][173] & ~x[36] & ~x[60] & ~x[62];
			partial_clause[9][174] 	= partial_clause_prev[9][174] & 1'b1;
			partial_clause[9][175] 	= partial_clause_prev[9][175] & 1'b1;
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & 1'b1;
			partial_clause[9][178] 	= partial_clause_prev[9][178] & 1'b1;
			partial_clause[9][179] 	= partial_clause_prev[9][179] & 1'b1;
			partial_clause[9][180] 	= partial_clause_prev[9][180] & 1'b1;
			partial_clause[9][181] 	= partial_clause_prev[9][181] & 1'b1;
			partial_clause[9][182] 	= partial_clause_prev[9][182] & 1'b1;
			partial_clause[9][183] 	= partial_clause_prev[9][183] & 1'b1;
			partial_clause[9][184] 	= partial_clause_prev[9][184] & ~x[9];
			partial_clause[9][185] 	= partial_clause_prev[9][185] & 1'b1;
			partial_clause[9][186] 	= partial_clause_prev[9][186] & 1'b1;
			partial_clause[9][187] 	= partial_clause_prev[9][187] & 1'b1;
			partial_clause[9][188] 	= partial_clause_prev[9][188] & 1'b1;
			partial_clause[9][189] 	= partial_clause_prev[9][189] & 1'b1;
			partial_clause[9][190] 	= partial_clause_prev[9][190] & 1'b1;
			partial_clause[9][191] 	= partial_clause_prev[9][191] & 1'b1;
			partial_clause[9][192] 	= partial_clause_prev[9][192] & x[1];
			partial_clause[9][193] 	= partial_clause_prev[9][193] & 1'b1;
			partial_clause[9][194] 	= partial_clause_prev[9][194] & x[1];
			partial_clause[9][195] 	= partial_clause_prev[9][195] & 1'b1;
			partial_clause[9][196] 	= partial_clause_prev[9][196] & 1'b1;
			partial_clause[9][197] 	= partial_clause_prev[9][197] & 1'b1;
			partial_clause[9][198] 	= partial_clause_prev[9][198] & 1'b1;
			partial_clause[9][199] 	= partial_clause_prev[9][199] & 1'b1;
		end
	end
endmodule


module HCB_5 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & ~x[31];
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & x[53];
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & ~x[57];
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & ~x[2] & ~x[58];
			partial_clause[0][11] 	= partial_clause_prev[0][11] & ~x[2];
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & x[37] & ~x[63];
			partial_clause[0][15] 	= partial_clause_prev[0][15] & ~x[59];
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & ~x[59];
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & x[34];
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & x[38];
			partial_clause[0][27] 	= partial_clause_prev[0][27] & ~x[60];
			partial_clause[0][28] 	= partial_clause_prev[0][28] & ~x[31];
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & x[11];
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & x[6];
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & x[27] & x[63];
			partial_clause[0][35] 	= partial_clause_prev[0][35] & x[53];
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & x[8];
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & x[35];
			partial_clause[0][49] 	= partial_clause_prev[0][49] & x[39];
			partial_clause[0][50] 	= partial_clause_prev[0][50] & ~x[60];
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & x[7];
			partial_clause[0][63] 	= partial_clause_prev[0][63] & ~x[30];
			partial_clause[0][64] 	= partial_clause_prev[0][64] & ~x[29];
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & x[33];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & ~x[58];
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & ~x[32];
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & x[63];
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & x[11];
			partial_clause[0][90] 	= partial_clause_prev[0][90] & x[28];
			partial_clause[0][91] 	= partial_clause_prev[0][91] & x[39];
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & x[53] & ~x[57];
			partial_clause[0][95] 	= partial_clause_prev[0][95] & x[50];
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & x[10];
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			partial_clause[0][100] 	= partial_clause_prev[0][100] & 1'b1;
			partial_clause[0][101] 	= partial_clause_prev[0][101] & ~x[31];
			partial_clause[0][102] 	= partial_clause_prev[0][102] & ~x[4] & ~x[27];
			partial_clause[0][103] 	= partial_clause_prev[0][103] & 1'b1;
			partial_clause[0][104] 	= partial_clause_prev[0][104] & ~x[11];
			partial_clause[0][105] 	= partial_clause_prev[0][105] & 1'b1;
			partial_clause[0][106] 	= partial_clause_prev[0][106] & 1'b1;
			partial_clause[0][107] 	= partial_clause_prev[0][107] & 1'b1;
			partial_clause[0][108] 	= partial_clause_prev[0][108] & ~x[30];
			partial_clause[0][109] 	= partial_clause_prev[0][109] & ~x[36];
			partial_clause[0][110] 	= partial_clause_prev[0][110] & ~x[49];
			partial_clause[0][111] 	= partial_clause_prev[0][111] & ~x[3];
			partial_clause[0][112] 	= partial_clause_prev[0][112] & ~x[35];
			partial_clause[0][113] 	= partial_clause_prev[0][113] & 1'b1;
			partial_clause[0][114] 	= partial_clause_prev[0][114] & 1'b1;
			partial_clause[0][115] 	= partial_clause_prev[0][115] & 1'b1;
			partial_clause[0][116] 	= partial_clause_prev[0][116] & 1'b1;
			partial_clause[0][117] 	= partial_clause_prev[0][117] & 1'b1;
			partial_clause[0][118] 	= partial_clause_prev[0][118] & 1'b1;
			partial_clause[0][119] 	= partial_clause_prev[0][119] & 1'b1;
			partial_clause[0][120] 	= partial_clause_prev[0][120] & 1'b1;
			partial_clause[0][121] 	= partial_clause_prev[0][121] & 1'b1;
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & 1'b1;
			partial_clause[0][124] 	= partial_clause_prev[0][124] & 1'b1;
			partial_clause[0][125] 	= partial_clause_prev[0][125] & 1'b1;
			partial_clause[0][126] 	= partial_clause_prev[0][126] & ~x[8] & x[58];
			partial_clause[0][127] 	= partial_clause_prev[0][127] & x[31];
			partial_clause[0][128] 	= partial_clause_prev[0][128] & 1'b1;
			partial_clause[0][129] 	= partial_clause_prev[0][129] & 1'b1;
			partial_clause[0][130] 	= partial_clause_prev[0][130] & 1'b1;
			partial_clause[0][131] 	= partial_clause_prev[0][131] & 1'b1;
			partial_clause[0][132] 	= partial_clause_prev[0][132] & 1'b1;
			partial_clause[0][133] 	= partial_clause_prev[0][133] & 1'b1;
			partial_clause[0][134] 	= partial_clause_prev[0][134] & 1'b1;
			partial_clause[0][135] 	= partial_clause_prev[0][135] & x[30];
			partial_clause[0][136] 	= partial_clause_prev[0][136] & 1'b1;
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & 1'b1;
			partial_clause[0][139] 	= partial_clause_prev[0][139] & x[4] & x[30];
			partial_clause[0][140] 	= partial_clause_prev[0][140] & 1'b1;
			partial_clause[0][141] 	= partial_clause_prev[0][141] & x[33];
			partial_clause[0][142] 	= partial_clause_prev[0][142] & 1'b1;
			partial_clause[0][143] 	= partial_clause_prev[0][143] & x[14];
			partial_clause[0][144] 	= partial_clause_prev[0][144] & 1'b1;
			partial_clause[0][145] 	= partial_clause_prev[0][145] & 1'b1;
			partial_clause[0][146] 	= partial_clause_prev[0][146] & ~x[3];
			partial_clause[0][147] 	= partial_clause_prev[0][147] & 1'b1;
			partial_clause[0][148] 	= partial_clause_prev[0][148] & 1'b1;
			partial_clause[0][149] 	= partial_clause_prev[0][149] & 1'b1;
			partial_clause[0][150] 	= partial_clause_prev[0][150] & ~x[4];
			partial_clause[0][151] 	= partial_clause_prev[0][151] & 1'b1;
			partial_clause[0][152] 	= partial_clause_prev[0][152] & 1'b1;
			partial_clause[0][153] 	= partial_clause_prev[0][153] & 1'b1;
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & 1'b1;
			partial_clause[0][156] 	= partial_clause_prev[0][156] & x[29];
			partial_clause[0][157] 	= partial_clause_prev[0][157] & 1'b1;
			partial_clause[0][158] 	= partial_clause_prev[0][158] & ~x[18];
			partial_clause[0][159] 	= partial_clause_prev[0][159] & 1'b1;
			partial_clause[0][160] 	= partial_clause_prev[0][160] & 1'b1;
			partial_clause[0][161] 	= partial_clause_prev[0][161] & 1'b1;
			partial_clause[0][162] 	= partial_clause_prev[0][162] & x[58] & x[59];
			partial_clause[0][163] 	= partial_clause_prev[0][163] & 1'b1;
			partial_clause[0][164] 	= partial_clause_prev[0][164] & x[4];
			partial_clause[0][165] 	= partial_clause_prev[0][165] & 1'b1;
			partial_clause[0][166] 	= partial_clause_prev[0][166] & 1'b1;
			partial_clause[0][167] 	= partial_clause_prev[0][167] & 1'b1;
			partial_clause[0][168] 	= partial_clause_prev[0][168] & 1'b1;
			partial_clause[0][169] 	= partial_clause_prev[0][169] & 1'b1;
			partial_clause[0][170] 	= partial_clause_prev[0][170] & x[60];
			partial_clause[0][171] 	= partial_clause_prev[0][171] & 1'b1;
			partial_clause[0][172] 	= partial_clause_prev[0][172] & 1'b1;
			partial_clause[0][173] 	= partial_clause_prev[0][173] & 1'b1;
			partial_clause[0][174] 	= partial_clause_prev[0][174] & ~x[25] & ~x[54] & ~x[55];
			partial_clause[0][175] 	= partial_clause_prev[0][175] & 1'b1;
			partial_clause[0][176] 	= partial_clause_prev[0][176] & 1'b1;
			partial_clause[0][177] 	= partial_clause_prev[0][177] & ~x[1];
			partial_clause[0][178] 	= partial_clause_prev[0][178] & 1'b1;
			partial_clause[0][179] 	= partial_clause_prev[0][179] & 1'b1;
			partial_clause[0][180] 	= partial_clause_prev[0][180] & x[59] & x[61];
			partial_clause[0][181] 	= partial_clause_prev[0][181] & 1'b1;
			partial_clause[0][182] 	= partial_clause_prev[0][182] & 1'b1;
			partial_clause[0][183] 	= partial_clause_prev[0][183] & 1'b1;
			partial_clause[0][184] 	= partial_clause_prev[0][184] & 1'b1;
			partial_clause[0][185] 	= partial_clause_prev[0][185] & 1'b1;
			partial_clause[0][186] 	= partial_clause_prev[0][186] & x[60];
			partial_clause[0][187] 	= partial_clause_prev[0][187] & 1'b1;
			partial_clause[0][188] 	= partial_clause_prev[0][188] & ~x[8] & ~x[34];
			partial_clause[0][189] 	= partial_clause_prev[0][189] & ~x[29] & ~x[39];
			partial_clause[0][190] 	= partial_clause_prev[0][190] & 1'b1;
			partial_clause[0][191] 	= partial_clause_prev[0][191] & 1'b1;
			partial_clause[0][192] 	= partial_clause_prev[0][192] & 1'b1;
			partial_clause[0][193] 	= partial_clause_prev[0][193] & 1'b1;
			partial_clause[0][194] 	= partial_clause_prev[0][194] & 1'b1;
			partial_clause[0][195] 	= partial_clause_prev[0][195] & 1'b1;
			partial_clause[0][196] 	= partial_clause_prev[0][196] & 1'b1;
			partial_clause[0][197] 	= partial_clause_prev[0][197] & ~x[9];
			partial_clause[0][198] 	= partial_clause_prev[0][198] & 1'b1;
			partial_clause[0][199] 	= partial_clause_prev[0][199] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[53];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & x[2] & ~x[35];
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & ~x[0] & x[3];
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & x[2];
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & x[30];
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & x[1];
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & ~x[61];
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & ~x[26] & ~x[28];
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & x[30];
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & ~x[5];
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & ~x[0];
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & x[4];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & x[1];
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & x[45];
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & x[59];
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & 1'b1;
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & x[31];
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & x[2] & x[3];
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & ~x[6];
			partial_clause[1][90] 	= partial_clause_prev[1][90] & ~x[27];
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			partial_clause[1][100] 	= partial_clause_prev[1][100] & 1'b1;
			partial_clause[1][101] 	= partial_clause_prev[1][101] & 1'b1;
			partial_clause[1][102] 	= partial_clause_prev[1][102] & ~x[31];
			partial_clause[1][103] 	= partial_clause_prev[1][103] & 1'b1;
			partial_clause[1][104] 	= partial_clause_prev[1][104] & 1'b1;
			partial_clause[1][105] 	= partial_clause_prev[1][105] & x[55];
			partial_clause[1][106] 	= partial_clause_prev[1][106] & 1'b1;
			partial_clause[1][107] 	= partial_clause_prev[1][107] & ~x[58];
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & 1'b1;
			partial_clause[1][110] 	= partial_clause_prev[1][110] & 1'b1;
			partial_clause[1][111] 	= partial_clause_prev[1][111] & 1'b1;
			partial_clause[1][112] 	= partial_clause_prev[1][112] & ~x[31];
			partial_clause[1][113] 	= partial_clause_prev[1][113] & 1'b1;
			partial_clause[1][114] 	= partial_clause_prev[1][114] & 1'b1;
			partial_clause[1][115] 	= partial_clause_prev[1][115] & 1'b1;
			partial_clause[1][116] 	= partial_clause_prev[1][116] & 1'b1;
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & 1'b1;
			partial_clause[1][119] 	= partial_clause_prev[1][119] & 1'b1;
			partial_clause[1][120] 	= partial_clause_prev[1][120] & 1'b1;
			partial_clause[1][121] 	= partial_clause_prev[1][121] & 1'b1;
			partial_clause[1][122] 	= partial_clause_prev[1][122] & 1'b1;
			partial_clause[1][123] 	= partial_clause_prev[1][123] & ~x[58];
			partial_clause[1][124] 	= partial_clause_prev[1][124] & 1'b1;
			partial_clause[1][125] 	= partial_clause_prev[1][125] & 1'b1;
			partial_clause[1][126] 	= partial_clause_prev[1][126] & 1'b1;
			partial_clause[1][127] 	= partial_clause_prev[1][127] & 1'b1;
			partial_clause[1][128] 	= partial_clause_prev[1][128] & 1'b1;
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & ~x[41];
			partial_clause[1][131] 	= partial_clause_prev[1][131] & 1'b1;
			partial_clause[1][132] 	= partial_clause_prev[1][132] & ~x[31];
			partial_clause[1][133] 	= partial_clause_prev[1][133] & 1'b1;
			partial_clause[1][134] 	= partial_clause_prev[1][134] & x[54];
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & x[54];
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & 1'b1;
			partial_clause[1][139] 	= partial_clause_prev[1][139] & 1'b1;
			partial_clause[1][140] 	= partial_clause_prev[1][140] & 1'b1;
			partial_clause[1][141] 	= partial_clause_prev[1][141] & 1'b1;
			partial_clause[1][142] 	= partial_clause_prev[1][142] & ~x[3];
			partial_clause[1][143] 	= partial_clause_prev[1][143] & 1'b1;
			partial_clause[1][144] 	= partial_clause_prev[1][144] & 1'b1;
			partial_clause[1][145] 	= partial_clause_prev[1][145] & ~x[3];
			partial_clause[1][146] 	= partial_clause_prev[1][146] & 1'b1;
			partial_clause[1][147] 	= partial_clause_prev[1][147] & 1'b1;
			partial_clause[1][148] 	= partial_clause_prev[1][148] & 1'b1;
			partial_clause[1][149] 	= partial_clause_prev[1][149] & 1'b1;
			partial_clause[1][150] 	= partial_clause_prev[1][150] & 1'b1;
			partial_clause[1][151] 	= partial_clause_prev[1][151] & 1'b1;
			partial_clause[1][152] 	= partial_clause_prev[1][152] & x[24];
			partial_clause[1][153] 	= partial_clause_prev[1][153] & 1'b1;
			partial_clause[1][154] 	= partial_clause_prev[1][154] & x[35];
			partial_clause[1][155] 	= partial_clause_prev[1][155] & 1'b1;
			partial_clause[1][156] 	= partial_clause_prev[1][156] & ~x[2];
			partial_clause[1][157] 	= partial_clause_prev[1][157] & 1'b1;
			partial_clause[1][158] 	= partial_clause_prev[1][158] & 1'b1;
			partial_clause[1][159] 	= partial_clause_prev[1][159] & x[27];
			partial_clause[1][160] 	= partial_clause_prev[1][160] & 1'b1;
			partial_clause[1][161] 	= partial_clause_prev[1][161] & 1'b1;
			partial_clause[1][162] 	= partial_clause_prev[1][162] & 1'b1;
			partial_clause[1][163] 	= partial_clause_prev[1][163] & 1'b1;
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & 1'b1;
			partial_clause[1][166] 	= partial_clause_prev[1][166] & 1'b1;
			partial_clause[1][167] 	= partial_clause_prev[1][167] & 1'b1;
			partial_clause[1][168] 	= partial_clause_prev[1][168] & ~x[3];
			partial_clause[1][169] 	= partial_clause_prev[1][169] & 1'b1;
			partial_clause[1][170] 	= partial_clause_prev[1][170] & 1'b1;
			partial_clause[1][171] 	= partial_clause_prev[1][171] & 1'b1;
			partial_clause[1][172] 	= partial_clause_prev[1][172] & 1'b1;
			partial_clause[1][173] 	= partial_clause_prev[1][173] & 1'b1;
			partial_clause[1][174] 	= partial_clause_prev[1][174] & 1'b1;
			partial_clause[1][175] 	= partial_clause_prev[1][175] & x[60];
			partial_clause[1][176] 	= partial_clause_prev[1][176] & 1'b1;
			partial_clause[1][177] 	= partial_clause_prev[1][177] & x[54];
			partial_clause[1][178] 	= partial_clause_prev[1][178] & 1'b1;
			partial_clause[1][179] 	= partial_clause_prev[1][179] & x[53];
			partial_clause[1][180] 	= partial_clause_prev[1][180] & 1'b1;
			partial_clause[1][181] 	= partial_clause_prev[1][181] & x[62];
			partial_clause[1][182] 	= partial_clause_prev[1][182] & 1'b1;
			partial_clause[1][183] 	= partial_clause_prev[1][183] & 1'b1;
			partial_clause[1][184] 	= partial_clause_prev[1][184] & ~x[58];
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & 1'b1;
			partial_clause[1][187] 	= partial_clause_prev[1][187] & 1'b1;
			partial_clause[1][188] 	= partial_clause_prev[1][188] & 1'b1;
			partial_clause[1][189] 	= partial_clause_prev[1][189] & 1'b1;
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & 1'b1;
			partial_clause[1][192] 	= partial_clause_prev[1][192] & ~x[30];
			partial_clause[1][193] 	= partial_clause_prev[1][193] & 1'b1;
			partial_clause[1][194] 	= partial_clause_prev[1][194] & 1'b1;
			partial_clause[1][195] 	= partial_clause_prev[1][195] & 1'b1;
			partial_clause[1][196] 	= partial_clause_prev[1][196] & 1'b1;
			partial_clause[1][197] 	= partial_clause_prev[1][197] & x[26];
			partial_clause[1][198] 	= partial_clause_prev[1][198] & 1'b1;
			partial_clause[1][199] 	= partial_clause_prev[1][199] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & ~x[2] & ~x[29] & ~x[56];
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & ~x[1];
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & ~x[1] & ~x[2] & ~x[31];
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & ~x[30];
			partial_clause[2][18] 	= partial_clause_prev[2][18] & ~x[28] & ~x[50];
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & ~x[30];
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & ~x[2];
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & ~x[2] & ~x[29] & ~x[53] & ~x[55];
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & ~x[54] & ~x[57];
			partial_clause[2][39] 	= partial_clause_prev[2][39] & ~x[1] & ~x[53];
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & ~x[0];
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & ~x[23];
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & ~x[22];
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & ~x[50];
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & 1'b1;
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & ~x[2];
			partial_clause[2][70] 	= partial_clause_prev[2][70] & ~x[29] & ~x[55] & ~x[57];
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & ~x[30] & ~x[56] & ~x[57];
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & ~x[22];
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & ~x[0] & ~x[2];
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & ~x[55];
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			partial_clause[2][100] 	= partial_clause_prev[2][100] & x[0] & ~x[24];
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & 1'b1;
			partial_clause[2][103] 	= partial_clause_prev[2][103] & x[23];
			partial_clause[2][104] 	= partial_clause_prev[2][104] & 1'b1;
			partial_clause[2][105] 	= partial_clause_prev[2][105] & 1'b1;
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & x[52];
			partial_clause[2][108] 	= partial_clause_prev[2][108] & 1'b1;
			partial_clause[2][109] 	= partial_clause_prev[2][109] & 1'b1;
			partial_clause[2][110] 	= partial_clause_prev[2][110] & 1'b1;
			partial_clause[2][111] 	= partial_clause_prev[2][111] & x[25];
			partial_clause[2][112] 	= partial_clause_prev[2][112] & x[55];
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & x[27];
			partial_clause[2][115] 	= partial_clause_prev[2][115] & x[18];
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & 1'b1;
			partial_clause[2][118] 	= partial_clause_prev[2][118] & 1'b1;
			partial_clause[2][119] 	= partial_clause_prev[2][119] & 1'b1;
			partial_clause[2][120] 	= partial_clause_prev[2][120] & 1'b1;
			partial_clause[2][121] 	= partial_clause_prev[2][121] & 1'b1;
			partial_clause[2][122] 	= partial_clause_prev[2][122] & 1'b1;
			partial_clause[2][123] 	= partial_clause_prev[2][123] & 1'b1;
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & 1'b1;
			partial_clause[2][126] 	= partial_clause_prev[2][126] & x[23];
			partial_clause[2][127] 	= partial_clause_prev[2][127] & x[53];
			partial_clause[2][128] 	= partial_clause_prev[2][128] & ~x[24] & x[27];
			partial_clause[2][129] 	= partial_clause_prev[2][129] & 1'b1;
			partial_clause[2][130] 	= partial_clause_prev[2][130] & 1'b1;
			partial_clause[2][131] 	= partial_clause_prev[2][131] & 1'b1;
			partial_clause[2][132] 	= partial_clause_prev[2][132] & 1'b1;
			partial_clause[2][133] 	= partial_clause_prev[2][133] & 1'b1;
			partial_clause[2][134] 	= partial_clause_prev[2][134] & 1'b1;
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & 1'b1;
			partial_clause[2][137] 	= partial_clause_prev[2][137] & 1'b1;
			partial_clause[2][138] 	= partial_clause_prev[2][138] & 1'b1;
			partial_clause[2][139] 	= partial_clause_prev[2][139] & 1'b1;
			partial_clause[2][140] 	= partial_clause_prev[2][140] & x[28];
			partial_clause[2][141] 	= partial_clause_prev[2][141] & ~x[23] & x[27];
			partial_clause[2][142] 	= partial_clause_prev[2][142] & 1'b1;
			partial_clause[2][143] 	= partial_clause_prev[2][143] & 1'b1;
			partial_clause[2][144] 	= partial_clause_prev[2][144] & x[49];
			partial_clause[2][145] 	= partial_clause_prev[2][145] & 1'b1;
			partial_clause[2][146] 	= partial_clause_prev[2][146] & x[54];
			partial_clause[2][147] 	= partial_clause_prev[2][147] & 1'b1;
			partial_clause[2][148] 	= partial_clause_prev[2][148] & 1'b1;
			partial_clause[2][149] 	= partial_clause_prev[2][149] & x[0];
			partial_clause[2][150] 	= partial_clause_prev[2][150] & 1'b1;
			partial_clause[2][151] 	= partial_clause_prev[2][151] & 1'b1;
			partial_clause[2][152] 	= partial_clause_prev[2][152] & x[50];
			partial_clause[2][153] 	= partial_clause_prev[2][153] & 1'b1;
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & x[29];
			partial_clause[2][156] 	= partial_clause_prev[2][156] & x[50];
			partial_clause[2][157] 	= partial_clause_prev[2][157] & x[53];
			partial_clause[2][158] 	= partial_clause_prev[2][158] & 1'b1;
			partial_clause[2][159] 	= partial_clause_prev[2][159] & 1'b1;
			partial_clause[2][160] 	= partial_clause_prev[2][160] & x[23];
			partial_clause[2][161] 	= partial_clause_prev[2][161] & 1'b1;
			partial_clause[2][162] 	= partial_clause_prev[2][162] & x[28];
			partial_clause[2][163] 	= partial_clause_prev[2][163] & 1'b1;
			partial_clause[2][164] 	= partial_clause_prev[2][164] & 1'b1;
			partial_clause[2][165] 	= partial_clause_prev[2][165] & 1'b1;
			partial_clause[2][166] 	= partial_clause_prev[2][166] & 1'b1;
			partial_clause[2][167] 	= partial_clause_prev[2][167] & 1'b1;
			partial_clause[2][168] 	= partial_clause_prev[2][168] & x[58];
			partial_clause[2][169] 	= partial_clause_prev[2][169] & 1'b1;
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & x[49];
			partial_clause[2][173] 	= partial_clause_prev[2][173] & 1'b1;
			partial_clause[2][174] 	= partial_clause_prev[2][174] & 1'b1;
			partial_clause[2][175] 	= partial_clause_prev[2][175] & 1'b1;
			partial_clause[2][176] 	= partial_clause_prev[2][176] & x[31];
			partial_clause[2][177] 	= partial_clause_prev[2][177] & 1'b1;
			partial_clause[2][178] 	= partial_clause_prev[2][178] & x[29];
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & 1'b1;
			partial_clause[2][181] 	= partial_clause_prev[2][181] & 1'b1;
			partial_clause[2][182] 	= partial_clause_prev[2][182] & x[55];
			partial_clause[2][183] 	= partial_clause_prev[2][183] & x[26] & ~x[50] & x[54];
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & 1'b1;
			partial_clause[2][186] 	= partial_clause_prev[2][186] & 1'b1;
			partial_clause[2][187] 	= partial_clause_prev[2][187] & 1'b1;
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & x[58];
			partial_clause[2][190] 	= partial_clause_prev[2][190] & 1'b1;
			partial_clause[2][191] 	= partial_clause_prev[2][191] & 1'b1;
			partial_clause[2][192] 	= partial_clause_prev[2][192] & x[24];
			partial_clause[2][193] 	= partial_clause_prev[2][193] & 1'b1;
			partial_clause[2][194] 	= partial_clause_prev[2][194] & 1'b1;
			partial_clause[2][195] 	= partial_clause_prev[2][195] & x[60];
			partial_clause[2][196] 	= partial_clause_prev[2][196] & 1'b1;
			partial_clause[2][197] 	= partial_clause_prev[2][197] & 1'b1;
			partial_clause[2][198] 	= partial_clause_prev[2][198] & 1'b1;
			partial_clause[2][199] 	= partial_clause_prev[2][199] & x[58] & x[59];
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & x[31] & x[56] & x[57] & x[58];
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & x[0] & x[1] & x[27];
			partial_clause[3][16] 	= partial_clause_prev[3][16] & x[0];
			partial_clause[3][17] 	= partial_clause_prev[3][17] & x[6];
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & x[6] & x[33];
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & x[2];
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & x[28];
			partial_clause[3][32] 	= partial_clause_prev[3][32] & x[42];
			partial_clause[3][33] 	= partial_clause_prev[3][33] & x[59];
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & ~x[24] & ~x[50];
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & ~x[51];
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & x[3] & x[56];
			partial_clause[3][42] 	= partial_clause_prev[3][42] & x[4];
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & x[5] & x[31] & x[58];
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & ~x[0] & ~x[23] & ~x[25];
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & x[59];
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & ~x[24];
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & x[13];
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & ~x[0] & ~x[25];
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & x[31];
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[40];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & ~x[25];
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & ~x[50];
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & x[28];
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & ~x[24];
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			partial_clause[3][100] 	= partial_clause_prev[3][100] & ~x[30];
			partial_clause[3][101] 	= partial_clause_prev[3][101] & x[50];
			partial_clause[3][102] 	= partial_clause_prev[3][102] & 1'b1;
			partial_clause[3][103] 	= partial_clause_prev[3][103] & 1'b1;
			partial_clause[3][104] 	= partial_clause_prev[3][104] & 1'b1;
			partial_clause[3][105] 	= partial_clause_prev[3][105] & 1'b1;
			partial_clause[3][106] 	= partial_clause_prev[3][106] & ~x[34];
			partial_clause[3][107] 	= partial_clause_prev[3][107] & 1'b1;
			partial_clause[3][108] 	= partial_clause_prev[3][108] & 1'b1;
			partial_clause[3][109] 	= partial_clause_prev[3][109] & 1'b1;
			partial_clause[3][110] 	= partial_clause_prev[3][110] & 1'b1;
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & 1'b1;
			partial_clause[3][113] 	= partial_clause_prev[3][113] & 1'b1;
			partial_clause[3][114] 	= partial_clause_prev[3][114] & 1'b1;
			partial_clause[3][115] 	= partial_clause_prev[3][115] & 1'b1;
			partial_clause[3][116] 	= partial_clause_prev[3][116] & 1'b1;
			partial_clause[3][117] 	= partial_clause_prev[3][117] & 1'b1;
			partial_clause[3][118] 	= partial_clause_prev[3][118] & 1'b1;
			partial_clause[3][119] 	= partial_clause_prev[3][119] & x[39];
			partial_clause[3][120] 	= partial_clause_prev[3][120] & x[24];
			partial_clause[3][121] 	= partial_clause_prev[3][121] & 1'b1;
			partial_clause[3][122] 	= partial_clause_prev[3][122] & ~x[2];
			partial_clause[3][123] 	= partial_clause_prev[3][123] & ~x[63];
			partial_clause[3][124] 	= partial_clause_prev[3][124] & 1'b1;
			partial_clause[3][125] 	= partial_clause_prev[3][125] & 1'b1;
			partial_clause[3][126] 	= partial_clause_prev[3][126] & ~x[3];
			partial_clause[3][127] 	= partial_clause_prev[3][127] & x[25];
			partial_clause[3][128] 	= partial_clause_prev[3][128] & ~x[5];
			partial_clause[3][129] 	= partial_clause_prev[3][129] & 1'b1;
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & 1'b1;
			partial_clause[3][132] 	= partial_clause_prev[3][132] & 1'b1;
			partial_clause[3][133] 	= partial_clause_prev[3][133] & 1'b1;
			partial_clause[3][134] 	= partial_clause_prev[3][134] & 1'b1;
			partial_clause[3][135] 	= partial_clause_prev[3][135] & 1'b1;
			partial_clause[3][136] 	= partial_clause_prev[3][136] & ~x[3] & ~x[59];
			partial_clause[3][137] 	= partial_clause_prev[3][137] & x[23];
			partial_clause[3][138] 	= partial_clause_prev[3][138] & 1'b1;
			partial_clause[3][139] 	= partial_clause_prev[3][139] & 1'b1;
			partial_clause[3][140] 	= partial_clause_prev[3][140] & 1'b1;
			partial_clause[3][141] 	= partial_clause_prev[3][141] & 1'b1;
			partial_clause[3][142] 	= partial_clause_prev[3][142] & 1'b1;
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & 1'b1;
			partial_clause[3][145] 	= partial_clause_prev[3][145] & 1'b1;
			partial_clause[3][146] 	= partial_clause_prev[3][146] & x[53];
			partial_clause[3][147] 	= partial_clause_prev[3][147] & ~x[30];
			partial_clause[3][148] 	= partial_clause_prev[3][148] & 1'b1;
			partial_clause[3][149] 	= partial_clause_prev[3][149] & 1'b1;
			partial_clause[3][150] 	= partial_clause_prev[3][150] & 1'b1;
			partial_clause[3][151] 	= partial_clause_prev[3][151] & ~x[5] & ~x[61];
			partial_clause[3][152] 	= partial_clause_prev[3][152] & 1'b1;
			partial_clause[3][153] 	= partial_clause_prev[3][153] & 1'b1;
			partial_clause[3][154] 	= partial_clause_prev[3][154] & x[23];
			partial_clause[3][155] 	= partial_clause_prev[3][155] & 1'b1;
			partial_clause[3][156] 	= partial_clause_prev[3][156] & 1'b1;
			partial_clause[3][157] 	= partial_clause_prev[3][157] & 1'b1;
			partial_clause[3][158] 	= partial_clause_prev[3][158] & ~x[32];
			partial_clause[3][159] 	= partial_clause_prev[3][159] & 1'b1;
			partial_clause[3][160] 	= partial_clause_prev[3][160] & 1'b1;
			partial_clause[3][161] 	= partial_clause_prev[3][161] & 1'b1;
			partial_clause[3][162] 	= partial_clause_prev[3][162] & 1'b1;
			partial_clause[3][163] 	= partial_clause_prev[3][163] & 1'b1;
			partial_clause[3][164] 	= partial_clause_prev[3][164] & 1'b1;
			partial_clause[3][165] 	= partial_clause_prev[3][165] & 1'b1;
			partial_clause[3][166] 	= partial_clause_prev[3][166] & 1'b1;
			partial_clause[3][167] 	= partial_clause_prev[3][167] & 1'b1;
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & x[51];
			partial_clause[3][170] 	= partial_clause_prev[3][170] & x[37];
			partial_clause[3][171] 	= partial_clause_prev[3][171] & 1'b1;
			partial_clause[3][172] 	= partial_clause_prev[3][172] & 1'b1;
			partial_clause[3][173] 	= partial_clause_prev[3][173] & 1'b1;
			partial_clause[3][174] 	= partial_clause_prev[3][174] & 1'b1;
			partial_clause[3][175] 	= partial_clause_prev[3][175] & 1'b1;
			partial_clause[3][176] 	= partial_clause_prev[3][176] & ~x[30];
			partial_clause[3][177] 	= partial_clause_prev[3][177] & x[27];
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & 1'b1;
			partial_clause[3][180] 	= partial_clause_prev[3][180] & 1'b1;
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & 1'b1;
			partial_clause[3][183] 	= partial_clause_prev[3][183] & 1'b1;
			partial_clause[3][184] 	= partial_clause_prev[3][184] & ~x[2] & ~x[58];
			partial_clause[3][185] 	= partial_clause_prev[3][185] & 1'b1;
			partial_clause[3][186] 	= partial_clause_prev[3][186] & x[27];
			partial_clause[3][187] 	= partial_clause_prev[3][187] & ~x[4] & ~x[60];
			partial_clause[3][188] 	= partial_clause_prev[3][188] & 1'b1;
			partial_clause[3][189] 	= partial_clause_prev[3][189] & 1'b1;
			partial_clause[3][190] 	= partial_clause_prev[3][190] & 1'b1;
			partial_clause[3][191] 	= partial_clause_prev[3][191] & ~x[25];
			partial_clause[3][192] 	= partial_clause_prev[3][192] & 1'b1;
			partial_clause[3][193] 	= partial_clause_prev[3][193] & 1'b1;
			partial_clause[3][194] 	= partial_clause_prev[3][194] & x[54];
			partial_clause[3][195] 	= partial_clause_prev[3][195] & 1'b1;
			partial_clause[3][196] 	= partial_clause_prev[3][196] & 1'b1;
			partial_clause[3][197] 	= partial_clause_prev[3][197] & 1'b1;
			partial_clause[3][198] 	= partial_clause_prev[3][198] & 1'b1;
			partial_clause[3][199] 	= partial_clause_prev[3][199] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & ~x[2];
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[2];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & ~x[2];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & x[45];
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & ~x[1];
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[1];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & ~x[1];
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & x[32] & ~x[35] & x[54];
			partial_clause[4][55] 	= partial_clause_prev[4][55] & ~x[1];
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & x[27] & x[32];
			partial_clause[4][65] 	= partial_clause_prev[4][65] & ~x[9];
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & ~x[39] & x[53];
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & x[25];
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & x[4];
			partial_clause[4][80] 	= partial_clause_prev[4][80] & ~x[30];
			partial_clause[4][81] 	= partial_clause_prev[4][81] & x[28];
			partial_clause[4][82] 	= partial_clause_prev[4][82] & ~x[2];
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & x[53];
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & x[54];
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & x[26] & x[53];
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			partial_clause[4][100] 	= partial_clause_prev[4][100] & 1'b1;
			partial_clause[4][101] 	= partial_clause_prev[4][101] & 1'b1;
			partial_clause[4][102] 	= partial_clause_prev[4][102] & 1'b1;
			partial_clause[4][103] 	= partial_clause_prev[4][103] & ~x[4];
			partial_clause[4][104] 	= partial_clause_prev[4][104] & 1'b1;
			partial_clause[4][105] 	= partial_clause_prev[4][105] & 1'b1;
			partial_clause[4][106] 	= partial_clause_prev[4][106] & 1'b1;
			partial_clause[4][107] 	= partial_clause_prev[4][107] & 1'b1;
			partial_clause[4][108] 	= partial_clause_prev[4][108] & ~x[55];
			partial_clause[4][109] 	= partial_clause_prev[4][109] & 1'b1;
			partial_clause[4][110] 	= partial_clause_prev[4][110] & ~x[26] & ~x[28] & ~x[49];
			partial_clause[4][111] 	= partial_clause_prev[4][111] & 1'b1;
			partial_clause[4][112] 	= partial_clause_prev[4][112] & 1'b1;
			partial_clause[4][113] 	= partial_clause_prev[4][113] & 1'b1;
			partial_clause[4][114] 	= partial_clause_prev[4][114] & 1'b1;
			partial_clause[4][115] 	= partial_clause_prev[4][115] & 1'b1;
			partial_clause[4][116] 	= partial_clause_prev[4][116] & 1'b1;
			partial_clause[4][117] 	= partial_clause_prev[4][117] & 1'b1;
			partial_clause[4][118] 	= partial_clause_prev[4][118] & 1'b1;
			partial_clause[4][119] 	= partial_clause_prev[4][119] & 1'b1;
			partial_clause[4][120] 	= partial_clause_prev[4][120] & ~x[52];
			partial_clause[4][121] 	= partial_clause_prev[4][121] & ~x[45] & ~x[55];
			partial_clause[4][122] 	= partial_clause_prev[4][122] & 1'b1;
			partial_clause[4][123] 	= partial_clause_prev[4][123] & 1'b1;
			partial_clause[4][124] 	= partial_clause_prev[4][124] & 1'b1;
			partial_clause[4][125] 	= partial_clause_prev[4][125] & 1'b1;
			partial_clause[4][126] 	= partial_clause_prev[4][126] & 1'b1;
			partial_clause[4][127] 	= partial_clause_prev[4][127] & 1'b1;
			partial_clause[4][128] 	= partial_clause_prev[4][128] & 1'b1;
			partial_clause[4][129] 	= partial_clause_prev[4][129] & 1'b1;
			partial_clause[4][130] 	= partial_clause_prev[4][130] & 1'b1;
			partial_clause[4][131] 	= partial_clause_prev[4][131] & ~x[0];
			partial_clause[4][132] 	= partial_clause_prev[4][132] & 1'b1;
			partial_clause[4][133] 	= partial_clause_prev[4][133] & ~x[23] & ~x[26] & ~x[27];
			partial_clause[4][134] 	= partial_clause_prev[4][134] & 1'b1;
			partial_clause[4][135] 	= partial_clause_prev[4][135] & 1'b1;
			partial_clause[4][136] 	= partial_clause_prev[4][136] & 1'b1;
			partial_clause[4][137] 	= partial_clause_prev[4][137] & ~x[53] & ~x[54];
			partial_clause[4][138] 	= partial_clause_prev[4][138] & ~x[61];
			partial_clause[4][139] 	= partial_clause_prev[4][139] & 1'b1;
			partial_clause[4][140] 	= partial_clause_prev[4][140] & 1'b1;
			partial_clause[4][141] 	= partial_clause_prev[4][141] & 1'b1;
			partial_clause[4][142] 	= partial_clause_prev[4][142] & 1'b1;
			partial_clause[4][143] 	= partial_clause_prev[4][143] & 1'b1;
			partial_clause[4][144] 	= partial_clause_prev[4][144] & 1'b1;
			partial_clause[4][145] 	= partial_clause_prev[4][145] & 1'b1;
			partial_clause[4][146] 	= partial_clause_prev[4][146] & 1'b1;
			partial_clause[4][147] 	= partial_clause_prev[4][147] & 1'b1;
			partial_clause[4][148] 	= partial_clause_prev[4][148] & 1'b1;
			partial_clause[4][149] 	= partial_clause_prev[4][149] & 1'b1;
			partial_clause[4][150] 	= partial_clause_prev[4][150] & ~x[56];
			partial_clause[4][151] 	= partial_clause_prev[4][151] & 1'b1;
			partial_clause[4][152] 	= partial_clause_prev[4][152] & 1'b1;
			partial_clause[4][153] 	= partial_clause_prev[4][153] & 1'b1;
			partial_clause[4][154] 	= partial_clause_prev[4][154] & 1'b1;
			partial_clause[4][155] 	= partial_clause_prev[4][155] & 1'b1;
			partial_clause[4][156] 	= partial_clause_prev[4][156] & 1'b1;
			partial_clause[4][157] 	= partial_clause_prev[4][157] & 1'b1;
			partial_clause[4][158] 	= partial_clause_prev[4][158] & 1'b1;
			partial_clause[4][159] 	= partial_clause_prev[4][159] & 1'b1;
			partial_clause[4][160] 	= partial_clause_prev[4][160] & 1'b1;
			partial_clause[4][161] 	= partial_clause_prev[4][161] & 1'b1;
			partial_clause[4][162] 	= partial_clause_prev[4][162] & 1'b1;
			partial_clause[4][163] 	= partial_clause_prev[4][163] & 1'b1;
			partial_clause[4][164] 	= partial_clause_prev[4][164] & 1'b1;
			partial_clause[4][165] 	= partial_clause_prev[4][165] & 1'b1;
			partial_clause[4][166] 	= partial_clause_prev[4][166] & 1'b1;
			partial_clause[4][167] 	= partial_clause_prev[4][167] & 1'b1;
			partial_clause[4][168] 	= partial_clause_prev[4][168] & 1'b1;
			partial_clause[4][169] 	= partial_clause_prev[4][169] & 1'b1;
			partial_clause[4][170] 	= partial_clause_prev[4][170] & ~x[60];
			partial_clause[4][171] 	= partial_clause_prev[4][171] & 1'b1;
			partial_clause[4][172] 	= partial_clause_prev[4][172] & 1'b1;
			partial_clause[4][173] 	= partial_clause_prev[4][173] & 1'b1;
			partial_clause[4][174] 	= partial_clause_prev[4][174] & 1'b1;
			partial_clause[4][175] 	= partial_clause_prev[4][175] & 1'b1;
			partial_clause[4][176] 	= partial_clause_prev[4][176] & 1'b1;
			partial_clause[4][177] 	= partial_clause_prev[4][177] & 1'b1;
			partial_clause[4][178] 	= partial_clause_prev[4][178] & 1'b1;
			partial_clause[4][179] 	= partial_clause_prev[4][179] & 1'b1;
			partial_clause[4][180] 	= partial_clause_prev[4][180] & ~x[54];
			partial_clause[4][181] 	= partial_clause_prev[4][181] & 1'b1;
			partial_clause[4][182] 	= partial_clause_prev[4][182] & 1'b1;
			partial_clause[4][183] 	= partial_clause_prev[4][183] & 1'b1;
			partial_clause[4][184] 	= partial_clause_prev[4][184] & 1'b1;
			partial_clause[4][185] 	= partial_clause_prev[4][185] & 1'b1;
			partial_clause[4][186] 	= partial_clause_prev[4][186] & ~x[61];
			partial_clause[4][187] 	= partial_clause_prev[4][187] & 1'b1;
			partial_clause[4][188] 	= partial_clause_prev[4][188] & 1'b1;
			partial_clause[4][189] 	= partial_clause_prev[4][189] & 1'b1;
			partial_clause[4][190] 	= partial_clause_prev[4][190] & ~x[0] & ~x[24] & ~x[25];
			partial_clause[4][191] 	= partial_clause_prev[4][191] & 1'b1;
			partial_clause[4][192] 	= partial_clause_prev[4][192] & 1'b1;
			partial_clause[4][193] 	= partial_clause_prev[4][193] & 1'b1;
			partial_clause[4][194] 	= partial_clause_prev[4][194] & 1'b1;
			partial_clause[4][195] 	= partial_clause_prev[4][195] & 1'b1;
			partial_clause[4][196] 	= partial_clause_prev[4][196] & 1'b1;
			partial_clause[4][197] 	= partial_clause_prev[4][197] & 1'b1;
			partial_clause[4][198] 	= partial_clause_prev[4][198] & 1'b1;
			partial_clause[4][199] 	= partial_clause_prev[4][199] & ~x[55];
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & x[4];
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & ~x[8] & ~x[39];
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & ~x[4] & ~x[34];
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & ~x[31];
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & ~x[9];
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & ~x[10];
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & ~x[9];
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & ~x[61] & ~x[62];
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & ~x[8];
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & ~x[60] & ~x[61];
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & ~x[37] & ~x[39];
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & ~x[8] & ~x[10] & ~x[11];
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & ~x[2] & ~x[3] & ~x[5];
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & x[1];
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & ~x[6] & ~x[7] & ~x[38];
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & ~x[61];
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & ~x[8];
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & ~x[10] & ~x[11];
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & ~x[11];
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			partial_clause[5][100] 	= partial_clause_prev[5][100] & 1'b1;
			partial_clause[5][101] 	= partial_clause_prev[5][101] & 1'b1;
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & 1'b1;
			partial_clause[5][104] 	= partial_clause_prev[5][104] & 1'b1;
			partial_clause[5][105] 	= partial_clause_prev[5][105] & x[9];
			partial_clause[5][106] 	= partial_clause_prev[5][106] & 1'b1;
			partial_clause[5][107] 	= partial_clause_prev[5][107] & 1'b1;
			partial_clause[5][108] 	= partial_clause_prev[5][108] & 1'b1;
			partial_clause[5][109] 	= partial_clause_prev[5][109] & ~x[36];
			partial_clause[5][110] 	= partial_clause_prev[5][110] & 1'b1;
			partial_clause[5][111] 	= partial_clause_prev[5][111] & 1'b1;
			partial_clause[5][112] 	= partial_clause_prev[5][112] & 1'b1;
			partial_clause[5][113] 	= partial_clause_prev[5][113] & 1'b1;
			partial_clause[5][114] 	= partial_clause_prev[5][114] & 1'b1;
			partial_clause[5][115] 	= partial_clause_prev[5][115] & x[38];
			partial_clause[5][116] 	= partial_clause_prev[5][116] & 1'b1;
			partial_clause[5][117] 	= partial_clause_prev[5][117] & 1'b1;
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & 1'b1;
			partial_clause[5][120] 	= partial_clause_prev[5][120] & x[38];
			partial_clause[5][121] 	= partial_clause_prev[5][121] & x[35];
			partial_clause[5][122] 	= partial_clause_prev[5][122] & 1'b1;
			partial_clause[5][123] 	= partial_clause_prev[5][123] & 1'b1;
			partial_clause[5][124] 	= partial_clause_prev[5][124] & 1'b1;
			partial_clause[5][125] 	= partial_clause_prev[5][125] & x[4] & x[59];
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & x[59];
			partial_clause[5][128] 	= partial_clause_prev[5][128] & 1'b1;
			partial_clause[5][129] 	= partial_clause_prev[5][129] & 1'b1;
			partial_clause[5][130] 	= partial_clause_prev[5][130] & ~x[4] & ~x[29] & ~x[56];
			partial_clause[5][131] 	= partial_clause_prev[5][131] & 1'b1;
			partial_clause[5][132] 	= partial_clause_prev[5][132] & 1'b1;
			partial_clause[5][133] 	= partial_clause_prev[5][133] & 1'b1;
			partial_clause[5][134] 	= partial_clause_prev[5][134] & 1'b1;
			partial_clause[5][135] 	= partial_clause_prev[5][135] & x[39];
			partial_clause[5][136] 	= partial_clause_prev[5][136] & x[8];
			partial_clause[5][137] 	= partial_clause_prev[5][137] & 1'b1;
			partial_clause[5][138] 	= partial_clause_prev[5][138] & 1'b1;
			partial_clause[5][139] 	= partial_clause_prev[5][139] & 1'b1;
			partial_clause[5][140] 	= partial_clause_prev[5][140] & ~x[3] & ~x[57];
			partial_clause[5][141] 	= partial_clause_prev[5][141] & 1'b1;
			partial_clause[5][142] 	= partial_clause_prev[5][142] & x[37];
			partial_clause[5][143] 	= partial_clause_prev[5][143] & 1'b1;
			partial_clause[5][144] 	= partial_clause_prev[5][144] & x[33];
			partial_clause[5][145] 	= partial_clause_prev[5][145] & 1'b1;
			partial_clause[5][146] 	= partial_clause_prev[5][146] & 1'b1;
			partial_clause[5][147] 	= partial_clause_prev[5][147] & x[4];
			partial_clause[5][148] 	= partial_clause_prev[5][148] & 1'b1;
			partial_clause[5][149] 	= partial_clause_prev[5][149] & 1'b1;
			partial_clause[5][150] 	= partial_clause_prev[5][150] & 1'b1;
			partial_clause[5][151] 	= partial_clause_prev[5][151] & x[62];
			partial_clause[5][152] 	= partial_clause_prev[5][152] & ~x[24];
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & 1'b1;
			partial_clause[5][155] 	= partial_clause_prev[5][155] & 1'b1;
			partial_clause[5][156] 	= partial_clause_prev[5][156] & x[35];
			partial_clause[5][157] 	= partial_clause_prev[5][157] & ~x[0];
			partial_clause[5][158] 	= partial_clause_prev[5][158] & 1'b1;
			partial_clause[5][159] 	= partial_clause_prev[5][159] & 1'b1;
			partial_clause[5][160] 	= partial_clause_prev[5][160] & 1'b1;
			partial_clause[5][161] 	= partial_clause_prev[5][161] & ~x[0] & ~x[28];
			partial_clause[5][162] 	= partial_clause_prev[5][162] & 1'b1;
			partial_clause[5][163] 	= partial_clause_prev[5][163] & x[39];
			partial_clause[5][164] 	= partial_clause_prev[5][164] & x[3];
			partial_clause[5][165] 	= partial_clause_prev[5][165] & 1'b1;
			partial_clause[5][166] 	= partial_clause_prev[5][166] & 1'b1;
			partial_clause[5][167] 	= partial_clause_prev[5][167] & 1'b1;
			partial_clause[5][168] 	= partial_clause_prev[5][168] & x[34];
			partial_clause[5][169] 	= partial_clause_prev[5][169] & 1'b1;
			partial_clause[5][170] 	= partial_clause_prev[5][170] & 1'b1;
			partial_clause[5][171] 	= partial_clause_prev[5][171] & 1'b1;
			partial_clause[5][172] 	= partial_clause_prev[5][172] & ~x[31];
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & x[8];
			partial_clause[5][175] 	= partial_clause_prev[5][175] & x[11];
			partial_clause[5][176] 	= partial_clause_prev[5][176] & 1'b1;
			partial_clause[5][177] 	= partial_clause_prev[5][177] & x[5];
			partial_clause[5][178] 	= partial_clause_prev[5][178] & 1'b1;
			partial_clause[5][179] 	= partial_clause_prev[5][179] & ~x[54];
			partial_clause[5][180] 	= partial_clause_prev[5][180] & ~x[12] & x[32] & ~x[50];
			partial_clause[5][181] 	= partial_clause_prev[5][181] & ~x[9];
			partial_clause[5][182] 	= partial_clause_prev[5][182] & x[7];
			partial_clause[5][183] 	= partial_clause_prev[5][183] & 1'b1;
			partial_clause[5][184] 	= partial_clause_prev[5][184] & 1'b1;
			partial_clause[5][185] 	= partial_clause_prev[5][185] & x[6];
			partial_clause[5][186] 	= partial_clause_prev[5][186] & 1'b1;
			partial_clause[5][187] 	= partial_clause_prev[5][187] & ~x[55];
			partial_clause[5][188] 	= partial_clause_prev[5][188] & x[38];
			partial_clause[5][189] 	= partial_clause_prev[5][189] & 1'b1;
			partial_clause[5][190] 	= partial_clause_prev[5][190] & ~x[0] & ~x[27];
			partial_clause[5][191] 	= partial_clause_prev[5][191] & 1'b1;
			partial_clause[5][192] 	= partial_clause_prev[5][192] & x[40];
			partial_clause[5][193] 	= partial_clause_prev[5][193] & 1'b1;
			partial_clause[5][194] 	= partial_clause_prev[5][194] & x[39];
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & 1'b1;
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & x[38];
			partial_clause[5][199] 	= partial_clause_prev[5][199] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & ~x[10];
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & x[55];
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & x[53];
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & x[1] & ~x[6] & ~x[10] & x[28];
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & ~x[3] & ~x[30];
			partial_clause[6][25] 	= partial_clause_prev[6][25] & x[7] & x[38];
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & x[1];
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & x[37];
			partial_clause[6][45] 	= partial_clause_prev[6][45] & ~x[4];
			partial_clause[6][46] 	= partial_clause_prev[6][46] & x[54];
			partial_clause[6][47] 	= partial_clause_prev[6][47] & x[1];
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & ~x[2];
			partial_clause[6][53] 	= partial_clause_prev[6][53] & ~x[4] & ~x[7];
			partial_clause[6][54] 	= partial_clause_prev[6][54] & ~x[38];
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & ~x[22] & x[27];
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & ~x[3] & ~x[4] & ~x[5] & ~x[7];
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & x[39];
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & x[55];
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & x[50];
			partial_clause[6][100] 	= partial_clause_prev[6][100] & 1'b1;
			partial_clause[6][101] 	= partial_clause_prev[6][101] & 1'b1;
			partial_clause[6][102] 	= partial_clause_prev[6][102] & 1'b1;
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & 1'b1;
			partial_clause[6][105] 	= partial_clause_prev[6][105] & 1'b1;
			partial_clause[6][106] 	= partial_clause_prev[6][106] & x[32] & ~x[36];
			partial_clause[6][107] 	= partial_clause_prev[6][107] & 1'b1;
			partial_clause[6][108] 	= partial_clause_prev[6][108] & 1'b1;
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & ~x[3];
			partial_clause[6][111] 	= partial_clause_prev[6][111] & 1'b1;
			partial_clause[6][112] 	= partial_clause_prev[6][112] & 1'b1;
			partial_clause[6][113] 	= partial_clause_prev[6][113] & 1'b1;
			partial_clause[6][114] 	= partial_clause_prev[6][114] & 1'b1;
			partial_clause[6][115] 	= partial_clause_prev[6][115] & 1'b1;
			partial_clause[6][116] 	= partial_clause_prev[6][116] & 1'b1;
			partial_clause[6][117] 	= partial_clause_prev[6][117] & 1'b1;
			partial_clause[6][118] 	= partial_clause_prev[6][118] & 1'b1;
			partial_clause[6][119] 	= partial_clause_prev[6][119] & 1'b1;
			partial_clause[6][120] 	= partial_clause_prev[6][120] & 1'b1;
			partial_clause[6][121] 	= partial_clause_prev[6][121] & ~x[52];
			partial_clause[6][122] 	= partial_clause_prev[6][122] & 1'b1;
			partial_clause[6][123] 	= partial_clause_prev[6][123] & 1'b1;
			partial_clause[6][124] 	= partial_clause_prev[6][124] & 1'b1;
			partial_clause[6][125] 	= partial_clause_prev[6][125] & x[58];
			partial_clause[6][126] 	= partial_clause_prev[6][126] & ~x[30] & ~x[57];
			partial_clause[6][127] 	= partial_clause_prev[6][127] & 1'b1;
			partial_clause[6][128] 	= partial_clause_prev[6][128] & 1'b1;
			partial_clause[6][129] 	= partial_clause_prev[6][129] & x[8] & ~x[30] & ~x[59];
			partial_clause[6][130] 	= partial_clause_prev[6][130] & x[35];
			partial_clause[6][131] 	= partial_clause_prev[6][131] & 1'b1;
			partial_clause[6][132] 	= partial_clause_prev[6][132] & 1'b1;
			partial_clause[6][133] 	= partial_clause_prev[6][133] & 1'b1;
			partial_clause[6][134] 	= partial_clause_prev[6][134] & ~x[32];
			partial_clause[6][135] 	= partial_clause_prev[6][135] & 1'b1;
			partial_clause[6][136] 	= partial_clause_prev[6][136] & 1'b1;
			partial_clause[6][137] 	= partial_clause_prev[6][137] & ~x[31];
			partial_clause[6][138] 	= partial_clause_prev[6][138] & ~x[59];
			partial_clause[6][139] 	= partial_clause_prev[6][139] & 1'b1;
			partial_clause[6][140] 	= partial_clause_prev[6][140] & ~x[10] & ~x[37];
			partial_clause[6][141] 	= partial_clause_prev[6][141] & 1'b1;
			partial_clause[6][142] 	= partial_clause_prev[6][142] & x[5];
			partial_clause[6][143] 	= partial_clause_prev[6][143] & 1'b1;
			partial_clause[6][144] 	= partial_clause_prev[6][144] & 1'b1;
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & ~x[3];
			partial_clause[6][147] 	= partial_clause_prev[6][147] & 1'b1;
			partial_clause[6][148] 	= partial_clause_prev[6][148] & 1'b1;
			partial_clause[6][149] 	= partial_clause_prev[6][149] & 1'b1;
			partial_clause[6][150] 	= partial_clause_prev[6][150] & 1'b1;
			partial_clause[6][151] 	= partial_clause_prev[6][151] & ~x[53];
			partial_clause[6][152] 	= partial_clause_prev[6][152] & 1'b1;
			partial_clause[6][153] 	= partial_clause_prev[6][153] & 1'b1;
			partial_clause[6][154] 	= partial_clause_prev[6][154] & ~x[37];
			partial_clause[6][155] 	= partial_clause_prev[6][155] & 1'b1;
			partial_clause[6][156] 	= partial_clause_prev[6][156] & 1'b1;
			partial_clause[6][157] 	= partial_clause_prev[6][157] & 1'b1;
			partial_clause[6][158] 	= partial_clause_prev[6][158] & 1'b1;
			partial_clause[6][159] 	= partial_clause_prev[6][159] & 1'b1;
			partial_clause[6][160] 	= partial_clause_prev[6][160] & 1'b1;
			partial_clause[6][161] 	= partial_clause_prev[6][161] & 1'b1;
			partial_clause[6][162] 	= partial_clause_prev[6][162] & 1'b1;
			partial_clause[6][163] 	= partial_clause_prev[6][163] & 1'b1;
			partial_clause[6][164] 	= partial_clause_prev[6][164] & 1'b1;
			partial_clause[6][165] 	= partial_clause_prev[6][165] & 1'b1;
			partial_clause[6][166] 	= partial_clause_prev[6][166] & ~x[4];
			partial_clause[6][167] 	= partial_clause_prev[6][167] & ~x[27];
			partial_clause[6][168] 	= partial_clause_prev[6][168] & 1'b1;
			partial_clause[6][169] 	= partial_clause_prev[6][169] & 1'b1;
			partial_clause[6][170] 	= partial_clause_prev[6][170] & 1'b1;
			partial_clause[6][171] 	= partial_clause_prev[6][171] & 1'b1;
			partial_clause[6][172] 	= partial_clause_prev[6][172] & 1'b1;
			partial_clause[6][173] 	= partial_clause_prev[6][173] & 1'b1;
			partial_clause[6][174] 	= partial_clause_prev[6][174] & 1'b1;
			partial_clause[6][175] 	= partial_clause_prev[6][175] & 1'b1;
			partial_clause[6][176] 	= partial_clause_prev[6][176] & ~x[28];
			partial_clause[6][177] 	= partial_clause_prev[6][177] & 1'b1;
			partial_clause[6][178] 	= partial_clause_prev[6][178] & ~x[4] & x[35];
			partial_clause[6][179] 	= partial_clause_prev[6][179] & 1'b1;
			partial_clause[6][180] 	= partial_clause_prev[6][180] & 1'b1;
			partial_clause[6][181] 	= partial_clause_prev[6][181] & 1'b1;
			partial_clause[6][182] 	= partial_clause_prev[6][182] & 1'b1;
			partial_clause[6][183] 	= partial_clause_prev[6][183] & 1'b1;
			partial_clause[6][184] 	= partial_clause_prev[6][184] & 1'b1;
			partial_clause[6][185] 	= partial_clause_prev[6][185] & 1'b1;
			partial_clause[6][186] 	= partial_clause_prev[6][186] & 1'b1;
			partial_clause[6][187] 	= partial_clause_prev[6][187] & 1'b1;
			partial_clause[6][188] 	= partial_clause_prev[6][188] & 1'b1;
			partial_clause[6][189] 	= partial_clause_prev[6][189] & 1'b1;
			partial_clause[6][190] 	= partial_clause_prev[6][190] & 1'b1;
			partial_clause[6][191] 	= partial_clause_prev[6][191] & 1'b1;
			partial_clause[6][192] 	= partial_clause_prev[6][192] & 1'b1;
			partial_clause[6][193] 	= partial_clause_prev[6][193] & 1'b1;
			partial_clause[6][194] 	= partial_clause_prev[6][194] & ~x[52] & ~x[54] & ~x[55] & ~x[56];
			partial_clause[6][195] 	= partial_clause_prev[6][195] & 1'b1;
			partial_clause[6][196] 	= partial_clause_prev[6][196] & ~x[52] & ~x[53];
			partial_clause[6][197] 	= partial_clause_prev[6][197] & 1'b1;
			partial_clause[6][198] 	= partial_clause_prev[6][198] & 1'b1;
			partial_clause[6][199] 	= partial_clause_prev[6][199] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & ~x[57];
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & ~x[30] & ~x[58];
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & ~x[57];
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & ~x[30];
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & ~x[59];
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & ~x[25];
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & ~x[23] & ~x[28] & ~x[54];
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & x[1];
			partial_clause[7][38] 	= partial_clause_prev[7][38] & ~x[27] & ~x[28] & ~x[53];
			partial_clause[7][39] 	= partial_clause_prev[7][39] & ~x[25] & ~x[27];
			partial_clause[7][40] 	= partial_clause_prev[7][40] & ~x[27] & x[32] & ~x[50] & ~x[52];
			partial_clause[7][41] 	= partial_clause_prev[7][41] & ~x[25];
			partial_clause[7][42] 	= partial_clause_prev[7][42] & ~x[25] & ~x[27] & ~x[51];
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & x[19];
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & x[47];
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & ~x[56] & ~x[58];
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & x[20];
			partial_clause[7][66] 	= partial_clause_prev[7][66] & x[20];
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & ~x[30];
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & ~x[30];
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & x[7];
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & x[19];
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & ~x[28];
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			partial_clause[7][100] 	= partial_clause_prev[7][100] & ~x[33];
			partial_clause[7][101] 	= partial_clause_prev[7][101] & 1'b1;
			partial_clause[7][102] 	= partial_clause_prev[7][102] & x[52];
			partial_clause[7][103] 	= partial_clause_prev[7][103] & 1'b1;
			partial_clause[7][104] 	= partial_clause_prev[7][104] & ~x[2];
			partial_clause[7][105] 	= partial_clause_prev[7][105] & ~x[1];
			partial_clause[7][106] 	= partial_clause_prev[7][106] & 1'b1;
			partial_clause[7][107] 	= partial_clause_prev[7][107] & 1'b1;
			partial_clause[7][108] 	= partial_clause_prev[7][108] & ~x[1];
			partial_clause[7][109] 	= partial_clause_prev[7][109] & ~x[35];
			partial_clause[7][110] 	= partial_clause_prev[7][110] & 1'b1;
			partial_clause[7][111] 	= partial_clause_prev[7][111] & 1'b1;
			partial_clause[7][112] 	= partial_clause_prev[7][112] & 1'b1;
			partial_clause[7][113] 	= partial_clause_prev[7][113] & ~x[5] & ~x[6];
			partial_clause[7][114] 	= partial_clause_prev[7][114] & 1'b1;
			partial_clause[7][115] 	= partial_clause_prev[7][115] & 1'b1;
			partial_clause[7][116] 	= partial_clause_prev[7][116] & 1'b1;
			partial_clause[7][117] 	= partial_clause_prev[7][117] & 1'b1;
			partial_clause[7][118] 	= partial_clause_prev[7][118] & 1'b1;
			partial_clause[7][119] 	= partial_clause_prev[7][119] & ~x[32];
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & x[24];
			partial_clause[7][123] 	= partial_clause_prev[7][123] & 1'b1;
			partial_clause[7][124] 	= partial_clause_prev[7][124] & 1'b1;
			partial_clause[7][125] 	= partial_clause_prev[7][125] & 1'b1;
			partial_clause[7][126] 	= partial_clause_prev[7][126] & 1'b1;
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & 1'b1;
			partial_clause[7][129] 	= partial_clause_prev[7][129] & 1'b1;
			partial_clause[7][130] 	= partial_clause_prev[7][130] & 1'b1;
			partial_clause[7][131] 	= partial_clause_prev[7][131] & 1'b1;
			partial_clause[7][132] 	= partial_clause_prev[7][132] & 1'b1;
			partial_clause[7][133] 	= partial_clause_prev[7][133] & 1'b1;
			partial_clause[7][134] 	= partial_clause_prev[7][134] & 1'b1;
			partial_clause[7][135] 	= partial_clause_prev[7][135] & ~x[9] & x[57];
			partial_clause[7][136] 	= partial_clause_prev[7][136] & 1'b1;
			partial_clause[7][137] 	= partial_clause_prev[7][137] & 1'b1;
			partial_clause[7][138] 	= partial_clause_prev[7][138] & 1'b1;
			partial_clause[7][139] 	= partial_clause_prev[7][139] & 1'b1;
			partial_clause[7][140] 	= partial_clause_prev[7][140] & 1'b1;
			partial_clause[7][141] 	= partial_clause_prev[7][141] & 1'b1;
			partial_clause[7][142] 	= partial_clause_prev[7][142] & x[25];
			partial_clause[7][143] 	= partial_clause_prev[7][143] & 1'b1;
			partial_clause[7][144] 	= partial_clause_prev[7][144] & 1'b1;
			partial_clause[7][145] 	= partial_clause_prev[7][145] & 1'b1;
			partial_clause[7][146] 	= partial_clause_prev[7][146] & 1'b1;
			partial_clause[7][147] 	= partial_clause_prev[7][147] & 1'b1;
			partial_clause[7][148] 	= partial_clause_prev[7][148] & 1'b1;
			partial_clause[7][149] 	= partial_clause_prev[7][149] & 1'b1;
			partial_clause[7][150] 	= partial_clause_prev[7][150] & ~x[2];
			partial_clause[7][151] 	= partial_clause_prev[7][151] & 1'b1;
			partial_clause[7][152] 	= partial_clause_prev[7][152] & 1'b1;
			partial_clause[7][153] 	= partial_clause_prev[7][153] & x[53];
			partial_clause[7][154] 	= partial_clause_prev[7][154] & 1'b1;
			partial_clause[7][155] 	= partial_clause_prev[7][155] & x[54];
			partial_clause[7][156] 	= partial_clause_prev[7][156] & 1'b1;
			partial_clause[7][157] 	= partial_clause_prev[7][157] & 1'b1;
			partial_clause[7][158] 	= partial_clause_prev[7][158] & 1'b1;
			partial_clause[7][159] 	= partial_clause_prev[7][159] & 1'b1;
			partial_clause[7][160] 	= partial_clause_prev[7][160] & 1'b1;
			partial_clause[7][161] 	= partial_clause_prev[7][161] & 1'b1;
			partial_clause[7][162] 	= partial_clause_prev[7][162] & 1'b1;
			partial_clause[7][163] 	= partial_clause_prev[7][163] & 1'b1;
			partial_clause[7][164] 	= partial_clause_prev[7][164] & 1'b1;
			partial_clause[7][165] 	= partial_clause_prev[7][165] & 1'b1;
			partial_clause[7][166] 	= partial_clause_prev[7][166] & x[30] & x[57];
			partial_clause[7][167] 	= partial_clause_prev[7][167] & 1'b1;
			partial_clause[7][168] 	= partial_clause_prev[7][168] & 1'b1;
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & x[55];
			partial_clause[7][171] 	= partial_clause_prev[7][171] & 1'b1;
			partial_clause[7][172] 	= partial_clause_prev[7][172] & 1'b1;
			partial_clause[7][173] 	= partial_clause_prev[7][173] & ~x[3];
			partial_clause[7][174] 	= partial_clause_prev[7][174] & 1'b1;
			partial_clause[7][175] 	= partial_clause_prev[7][175] & 1'b1;
			partial_clause[7][176] 	= partial_clause_prev[7][176] & 1'b1;
			partial_clause[7][177] 	= partial_clause_prev[7][177] & 1'b1;
			partial_clause[7][178] 	= partial_clause_prev[7][178] & ~x[8] & x[29] & ~x[50];
			partial_clause[7][179] 	= partial_clause_prev[7][179] & 1'b1;
			partial_clause[7][180] 	= partial_clause_prev[7][180] & x[52];
			partial_clause[7][181] 	= partial_clause_prev[7][181] & 1'b1;
			partial_clause[7][182] 	= partial_clause_prev[7][182] & 1'b1;
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & 1'b1;
			partial_clause[7][185] 	= partial_clause_prev[7][185] & ~x[38] & x[56];
			partial_clause[7][186] 	= partial_clause_prev[7][186] & ~x[4];
			partial_clause[7][187] 	= partial_clause_prev[7][187] & 1'b1;
			partial_clause[7][188] 	= partial_clause_prev[7][188] & x[25];
			partial_clause[7][189] 	= partial_clause_prev[7][189] & 1'b1;
			partial_clause[7][190] 	= partial_clause_prev[7][190] & ~x[21] & x[57];
			partial_clause[7][191] 	= partial_clause_prev[7][191] & 1'b1;
			partial_clause[7][192] 	= partial_clause_prev[7][192] & x[39];
			partial_clause[7][193] 	= partial_clause_prev[7][193] & 1'b1;
			partial_clause[7][194] 	= partial_clause_prev[7][194] & 1'b1;
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & ~x[21] & x[57];
			partial_clause[7][197] 	= partial_clause_prev[7][197] & 1'b1;
			partial_clause[7][198] 	= partial_clause_prev[7][198] & ~x[24];
			partial_clause[7][199] 	= partial_clause_prev[7][199] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & x[27];
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & x[30];
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & x[6];
			partial_clause[8][19] 	= partial_clause_prev[8][19] & x[35];
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & x[1] & x[30];
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & x[56];
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & x[10];
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & x[12];
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & x[7];
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & x[6] & ~x[53];
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & x[57];
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & x[9] & x[61];
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & x[37];
			partial_clause[8][64] 	= partial_clause_prev[8][64] & x[16];
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & x[11];
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & x[28] & ~x[53];
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & x[19];
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & x[58];
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & x[33] & ~x[54];
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & x[16];
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			partial_clause[8][100] 	= partial_clause_prev[8][100] & 1'b1;
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & 1'b1;
			partial_clause[8][103] 	= partial_clause_prev[8][103] & 1'b1;
			partial_clause[8][104] 	= partial_clause_prev[8][104] & x[17];
			partial_clause[8][105] 	= partial_clause_prev[8][105] & 1'b1;
			partial_clause[8][106] 	= partial_clause_prev[8][106] & 1'b1;
			partial_clause[8][107] 	= partial_clause_prev[8][107] & ~x[2] & ~x[20] & ~x[29] & ~x[56];
			partial_clause[8][108] 	= partial_clause_prev[8][108] & 1'b1;
			partial_clause[8][109] 	= partial_clause_prev[8][109] & 1'b1;
			partial_clause[8][110] 	= partial_clause_prev[8][110] & 1'b1;
			partial_clause[8][111] 	= partial_clause_prev[8][111] & 1'b1;
			partial_clause[8][112] 	= partial_clause_prev[8][112] & ~x[29] & ~x[56];
			partial_clause[8][113] 	= partial_clause_prev[8][113] & 1'b1;
			partial_clause[8][114] 	= partial_clause_prev[8][114] & ~x[11];
			partial_clause[8][115] 	= partial_clause_prev[8][115] & 1'b1;
			partial_clause[8][116] 	= partial_clause_prev[8][116] & 1'b1;
			partial_clause[8][117] 	= partial_clause_prev[8][117] & 1'b1;
			partial_clause[8][118] 	= partial_clause_prev[8][118] & 1'b1;
			partial_clause[8][119] 	= partial_clause_prev[8][119] & 1'b1;
			partial_clause[8][120] 	= partial_clause_prev[8][120] & 1'b1;
			partial_clause[8][121] 	= partial_clause_prev[8][121] & 1'b1;
			partial_clause[8][122] 	= partial_clause_prev[8][122] & 1'b1;
			partial_clause[8][123] 	= partial_clause_prev[8][123] & 1'b1;
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & 1'b1;
			partial_clause[8][126] 	= partial_clause_prev[8][126] & 1'b1;
			partial_clause[8][127] 	= partial_clause_prev[8][127] & 1'b1;
			partial_clause[8][128] 	= partial_clause_prev[8][128] & 1'b1;
			partial_clause[8][129] 	= partial_clause_prev[8][129] & 1'b1;
			partial_clause[8][130] 	= partial_clause_prev[8][130] & 1'b1;
			partial_clause[8][131] 	= partial_clause_prev[8][131] & 1'b1;
			partial_clause[8][132] 	= partial_clause_prev[8][132] & 1'b1;
			partial_clause[8][133] 	= partial_clause_prev[8][133] & ~x[25] & ~x[51];
			partial_clause[8][134] 	= partial_clause_prev[8][134] & 1'b1;
			partial_clause[8][135] 	= partial_clause_prev[8][135] & 1'b1;
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & ~x[58];
			partial_clause[8][138] 	= partial_clause_prev[8][138] & 1'b1;
			partial_clause[8][139] 	= partial_clause_prev[8][139] & 1'b1;
			partial_clause[8][140] 	= partial_clause_prev[8][140] & 1'b1;
			partial_clause[8][141] 	= partial_clause_prev[8][141] & 1'b1;
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & 1'b1;
			partial_clause[8][144] 	= partial_clause_prev[8][144] & 1'b1;
			partial_clause[8][145] 	= partial_clause_prev[8][145] & ~x[35];
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & 1'b1;
			partial_clause[8][148] 	= partial_clause_prev[8][148] & 1'b1;
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & 1'b1;
			partial_clause[8][151] 	= partial_clause_prev[8][151] & 1'b1;
			partial_clause[8][152] 	= partial_clause_prev[8][152] & 1'b1;
			partial_clause[8][153] 	= partial_clause_prev[8][153] & ~x[1] & ~x[28] & ~x[56];
			partial_clause[8][154] 	= partial_clause_prev[8][154] & 1'b1;
			partial_clause[8][155] 	= partial_clause_prev[8][155] & 1'b1;
			partial_clause[8][156] 	= partial_clause_prev[8][156] & ~x[30];
			partial_clause[8][157] 	= partial_clause_prev[8][157] & 1'b1;
			partial_clause[8][158] 	= partial_clause_prev[8][158] & 1'b1;
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & 1'b1;
			partial_clause[8][161] 	= partial_clause_prev[8][161] & 1'b1;
			partial_clause[8][162] 	= partial_clause_prev[8][162] & ~x[30];
			partial_clause[8][163] 	= partial_clause_prev[8][163] & ~x[29] & ~x[56];
			partial_clause[8][164] 	= partial_clause_prev[8][164] & ~x[0] & ~x[27] & ~x[55];
			partial_clause[8][165] 	= partial_clause_prev[8][165] & ~x[12];
			partial_clause[8][166] 	= partial_clause_prev[8][166] & 1'b1;
			partial_clause[8][167] 	= partial_clause_prev[8][167] & 1'b1;
			partial_clause[8][168] 	= partial_clause_prev[8][168] & 1'b1;
			partial_clause[8][169] 	= partial_clause_prev[8][169] & ~x[51];
			partial_clause[8][170] 	= partial_clause_prev[8][170] & 1'b1;
			partial_clause[8][171] 	= partial_clause_prev[8][171] & 1'b1;
			partial_clause[8][172] 	= partial_clause_prev[8][172] & 1'b1;
			partial_clause[8][173] 	= partial_clause_prev[8][173] & 1'b1;
			partial_clause[8][174] 	= partial_clause_prev[8][174] & 1'b1;
			partial_clause[8][175] 	= partial_clause_prev[8][175] & 1'b1;
			partial_clause[8][176] 	= partial_clause_prev[8][176] & 1'b1;
			partial_clause[8][177] 	= partial_clause_prev[8][177] & ~x[58];
			partial_clause[8][178] 	= partial_clause_prev[8][178] & 1'b1;
			partial_clause[8][179] 	= partial_clause_prev[8][179] & 1'b1;
			partial_clause[8][180] 	= partial_clause_prev[8][180] & 1'b1;
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & ~x[23] & ~x[37];
			partial_clause[8][183] 	= partial_clause_prev[8][183] & 1'b1;
			partial_clause[8][184] 	= partial_clause_prev[8][184] & 1'b1;
			partial_clause[8][185] 	= partial_clause_prev[8][185] & 1'b1;
			partial_clause[8][186] 	= partial_clause_prev[8][186] & ~x[59];
			partial_clause[8][187] 	= partial_clause_prev[8][187] & 1'b1;
			partial_clause[8][188] 	= partial_clause_prev[8][188] & ~x[60];
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & 1'b1;
			partial_clause[8][191] 	= partial_clause_prev[8][191] & 1'b1;
			partial_clause[8][192] 	= partial_clause_prev[8][192] & ~x[28];
			partial_clause[8][193] 	= partial_clause_prev[8][193] & 1'b1;
			partial_clause[8][194] 	= partial_clause_prev[8][194] & 1'b1;
			partial_clause[8][195] 	= partial_clause_prev[8][195] & 1'b1;
			partial_clause[8][196] 	= partial_clause_prev[8][196] & 1'b1;
			partial_clause[8][197] 	= partial_clause_prev[8][197] & 1'b1;
			partial_clause[8][198] 	= partial_clause_prev[8][198] & 1'b1;
			partial_clause[8][199] 	= partial_clause_prev[8][199] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & x[63];
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & x[21];
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & x[59];
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & x[49];
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & ~x[0];
			partial_clause[9][30] 	= partial_clause_prev[9][30] & ~x[1] & x[25];
			partial_clause[9][31] 	= partial_clause_prev[9][31] & x[52];
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & x[34];
			partial_clause[9][35] 	= partial_clause_prev[9][35] & 1'b1;
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & x[43];
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & x[16];
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & x[59];
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & x[34];
			partial_clause[9][71] 	= partial_clause_prev[9][71] & x[22];
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & x[21];
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & x[63];
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & ~x[28];
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
			partial_clause[9][100] 	= partial_clause_prev[9][100] & ~x[50] & ~x[60];
			partial_clause[9][101] 	= partial_clause_prev[9][101] & 1'b1;
			partial_clause[9][102] 	= partial_clause_prev[9][102] & 1'b1;
			partial_clause[9][103] 	= partial_clause_prev[9][103] & 1'b1;
			partial_clause[9][104] 	= partial_clause_prev[9][104] & 1'b1;
			partial_clause[9][105] 	= partial_clause_prev[9][105] & 1'b1;
			partial_clause[9][106] 	= partial_clause_prev[9][106] & 1'b1;
			partial_clause[9][107] 	= partial_clause_prev[9][107] & ~x[35];
			partial_clause[9][108] 	= partial_clause_prev[9][108] & 1'b1;
			partial_clause[9][109] 	= partial_clause_prev[9][109] & 1'b1;
			partial_clause[9][110] 	= partial_clause_prev[9][110] & 1'b1;
			partial_clause[9][111] 	= partial_clause_prev[9][111] & ~x[25] & ~x[50] & ~x[51];
			partial_clause[9][112] 	= partial_clause_prev[9][112] & 1'b1;
			partial_clause[9][113] 	= partial_clause_prev[9][113] & ~x[3];
			partial_clause[9][114] 	= partial_clause_prev[9][114] & 1'b1;
			partial_clause[9][115] 	= partial_clause_prev[9][115] & 1'b1;
			partial_clause[9][116] 	= partial_clause_prev[9][116] & ~x[60];
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & ~x[30];
			partial_clause[9][119] 	= partial_clause_prev[9][119] & ~x[22] & ~x[23];
			partial_clause[9][120] 	= partial_clause_prev[9][120] & 1'b1;
			partial_clause[9][121] 	= partial_clause_prev[9][121] & 1'b1;
			partial_clause[9][122] 	= partial_clause_prev[9][122] & ~x[22] & ~x[23] & ~x[34] & ~x[35] & ~x[36];
			partial_clause[9][123] 	= partial_clause_prev[9][123] & 1'b1;
			partial_clause[9][124] 	= partial_clause_prev[9][124] & 1'b1;
			partial_clause[9][125] 	= partial_clause_prev[9][125] & ~x[0] & ~x[22] & ~x[24] & ~x[26];
			partial_clause[9][126] 	= partial_clause_prev[9][126] & 1'b1;
			partial_clause[9][127] 	= partial_clause_prev[9][127] & 1'b1;
			partial_clause[9][128] 	= partial_clause_prev[9][128] & 1'b1;
			partial_clause[9][129] 	= partial_clause_prev[9][129] & ~x[30];
			partial_clause[9][130] 	= partial_clause_prev[9][130] & 1'b1;
			partial_clause[9][131] 	= partial_clause_prev[9][131] & 1'b1;
			partial_clause[9][132] 	= partial_clause_prev[9][132] & ~x[7] & ~x[33] & ~x[36];
			partial_clause[9][133] 	= partial_clause_prev[9][133] & 1'b1;
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & 1'b1;
			partial_clause[9][138] 	= partial_clause_prev[9][138] & 1'b1;
			partial_clause[9][139] 	= partial_clause_prev[9][139] & 1'b1;
			partial_clause[9][140] 	= partial_clause_prev[9][140] & 1'b1;
			partial_clause[9][141] 	= partial_clause_prev[9][141] & 1'b1;
			partial_clause[9][142] 	= partial_clause_prev[9][142] & 1'b1;
			partial_clause[9][143] 	= partial_clause_prev[9][143] & 1'b1;
			partial_clause[9][144] 	= partial_clause_prev[9][144] & 1'b1;
			partial_clause[9][145] 	= partial_clause_prev[9][145] & 1'b1;
			partial_clause[9][146] 	= partial_clause_prev[9][146] & 1'b1;
			partial_clause[9][147] 	= partial_clause_prev[9][147] & ~x[23] & ~x[24];
			partial_clause[9][148] 	= partial_clause_prev[9][148] & ~x[29];
			partial_clause[9][149] 	= partial_clause_prev[9][149] & ~x[55];
			partial_clause[9][150] 	= partial_clause_prev[9][150] & 1'b1;
			partial_clause[9][151] 	= partial_clause_prev[9][151] & ~x[62];
			partial_clause[9][152] 	= partial_clause_prev[9][152] & 1'b1;
			partial_clause[9][153] 	= partial_clause_prev[9][153] & 1'b1;
			partial_clause[9][154] 	= partial_clause_prev[9][154] & ~x[51] & ~x[53] & ~x[54];
			partial_clause[9][155] 	= partial_clause_prev[9][155] & 1'b1;
			partial_clause[9][156] 	= partial_clause_prev[9][156] & 1'b1;
			partial_clause[9][157] 	= partial_clause_prev[9][157] & ~x[33] & ~x[34];
			partial_clause[9][158] 	= partial_clause_prev[9][158] & ~x[27] & ~x[53] & ~x[54];
			partial_clause[9][159] 	= partial_clause_prev[9][159] & 1'b1;
			partial_clause[9][160] 	= partial_clause_prev[9][160] & 1'b1;
			partial_clause[9][161] 	= partial_clause_prev[9][161] & 1'b1;
			partial_clause[9][162] 	= partial_clause_prev[9][162] & 1'b1;
			partial_clause[9][163] 	= partial_clause_prev[9][163] & 1'b1;
			partial_clause[9][164] 	= partial_clause_prev[9][164] & 1'b1;
			partial_clause[9][165] 	= partial_clause_prev[9][165] & ~x[22];
			partial_clause[9][166] 	= partial_clause_prev[9][166] & 1'b1;
			partial_clause[9][167] 	= partial_clause_prev[9][167] & 1'b1;
			partial_clause[9][168] 	= partial_clause_prev[9][168] & ~x[20];
			partial_clause[9][169] 	= partial_clause_prev[9][169] & 1'b1;
			partial_clause[9][170] 	= partial_clause_prev[9][170] & 1'b1;
			partial_clause[9][171] 	= partial_clause_prev[9][171] & 1'b1;
			partial_clause[9][172] 	= partial_clause_prev[9][172] & ~x[28] & ~x[54];
			partial_clause[9][173] 	= partial_clause_prev[9][173] & ~x[49];
			partial_clause[9][174] 	= partial_clause_prev[9][174] & 1'b1;
			partial_clause[9][175] 	= partial_clause_prev[9][175] & 1'b1;
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & 1'b1;
			partial_clause[9][178] 	= partial_clause_prev[9][178] & 1'b1;
			partial_clause[9][179] 	= partial_clause_prev[9][179] & 1'b1;
			partial_clause[9][180] 	= partial_clause_prev[9][180] & 1'b1;
			partial_clause[9][181] 	= partial_clause_prev[9][181] & 1'b1;
			partial_clause[9][182] 	= partial_clause_prev[9][182] & ~x[28] & ~x[55];
			partial_clause[9][183] 	= partial_clause_prev[9][183] & 1'b1;
			partial_clause[9][184] 	= partial_clause_prev[9][184] & 1'b1;
			partial_clause[9][185] 	= partial_clause_prev[9][185] & 1'b1;
			partial_clause[9][186] 	= partial_clause_prev[9][186] & 1'b1;
			partial_clause[9][187] 	= partial_clause_prev[9][187] & ~x[58];
			partial_clause[9][188] 	= partial_clause_prev[9][188] & 1'b1;
			partial_clause[9][189] 	= partial_clause_prev[9][189] & 1'b1;
			partial_clause[9][190] 	= partial_clause_prev[9][190] & 1'b1;
			partial_clause[9][191] 	= partial_clause_prev[9][191] & 1'b1;
			partial_clause[9][192] 	= partial_clause_prev[9][192] & 1'b1;
			partial_clause[9][193] 	= partial_clause_prev[9][193] & 1'b1;
			partial_clause[9][194] 	= partial_clause_prev[9][194] & 1'b1;
			partial_clause[9][195] 	= partial_clause_prev[9][195] & 1'b1;
			partial_clause[9][196] 	= partial_clause_prev[9][196] & ~x[32];
			partial_clause[9][197] 	= partial_clause_prev[9][197] & 1'b1;
			partial_clause[9][198] 	= partial_clause_prev[9][198] & 1'b1;
			partial_clause[9][199] 	= partial_clause_prev[9][199] & 1'b1;
		end
	end
endmodule


module HCB_6 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & x[30];
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & x[1];
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & ~x[21] & ~x[51];
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & ~x[50];
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & ~x[49];
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & x[1];
			partial_clause[0][22] 	= partial_clause_prev[0][22] & x[41];
			partial_clause[0][23] 	= partial_clause_prev[0][23] & x[46];
			partial_clause[0][24] 	= partial_clause_prev[0][24] & x[44];
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & ~x[47];
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & ~x[51];
			partial_clause[0][29] 	= partial_clause_prev[0][29] & x[60];
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & x[45];
			partial_clause[0][35] 	= partial_clause_prev[0][35] & ~x[25];
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & ~x[21] & ~x[50];
			partial_clause[0][47] 	= partial_clause_prev[0][47] & x[40];
			partial_clause[0][48] 	= partial_clause_prev[0][48] & x[45];
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & x[60];
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & x[18];
			partial_clause[0][54] 	= partial_clause_prev[0][54] & x[8];
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & x[4];
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & ~x[54];
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & x[18];
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & ~x[21] & ~x[25];
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & x[46];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & x[5];
			partial_clause[0][78] 	= partial_clause_prev[0][78] & x[16] & ~x[26];
			partial_clause[0][79] 	= partial_clause_prev[0][79] & x[6];
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & x[2];
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & ~x[26] & x[43];
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & x[27] & x[45];
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & ~x[26];
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & x[0];
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & x[43];
			partial_clause[0][99] 	= partial_clause_prev[0][99] & x[3];
			partial_clause[0][100] 	= partial_clause_prev[0][100] & 1'b1;
			partial_clause[0][101] 	= partial_clause_prev[0][101] & 1'b1;
			partial_clause[0][102] 	= partial_clause_prev[0][102] & 1'b1;
			partial_clause[0][103] 	= partial_clause_prev[0][103] & 1'b1;
			partial_clause[0][104] 	= partial_clause_prev[0][104] & 1'b1;
			partial_clause[0][105] 	= partial_clause_prev[0][105] & ~x[31];
			partial_clause[0][106] 	= partial_clause_prev[0][106] & 1'b1;
			partial_clause[0][107] 	= partial_clause_prev[0][107] & x[22];
			partial_clause[0][108] 	= partial_clause_prev[0][108] & ~x[31];
			partial_clause[0][109] 	= partial_clause_prev[0][109] & ~x[26] & ~x[30];
			partial_clause[0][110] 	= partial_clause_prev[0][110] & 1'b1;
			partial_clause[0][111] 	= partial_clause_prev[0][111] & 1'b1;
			partial_clause[0][112] 	= partial_clause_prev[0][112] & ~x[2] & ~x[3];
			partial_clause[0][113] 	= partial_clause_prev[0][113] & 1'b1;
			partial_clause[0][114] 	= partial_clause_prev[0][114] & x[22];
			partial_clause[0][115] 	= partial_clause_prev[0][115] & 1'b1;
			partial_clause[0][116] 	= partial_clause_prev[0][116] & 1'b1;
			partial_clause[0][117] 	= partial_clause_prev[0][117] & 1'b1;
			partial_clause[0][118] 	= partial_clause_prev[0][118] & 1'b1;
			partial_clause[0][119] 	= partial_clause_prev[0][119] & 1'b1;
			partial_clause[0][120] 	= partial_clause_prev[0][120] & x[23];
			partial_clause[0][121] 	= partial_clause_prev[0][121] & 1'b1;
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & ~x[46] & ~x[47];
			partial_clause[0][124] 	= partial_clause_prev[0][124] & 1'b1;
			partial_clause[0][125] 	= partial_clause_prev[0][125] & 1'b1;
			partial_clause[0][126] 	= partial_clause_prev[0][126] & 1'b1;
			partial_clause[0][127] 	= partial_clause_prev[0][127] & 1'b1;
			partial_clause[0][128] 	= partial_clause_prev[0][128] & 1'b1;
			partial_clause[0][129] 	= partial_clause_prev[0][129] & x[51];
			partial_clause[0][130] 	= partial_clause_prev[0][130] & 1'b1;
			partial_clause[0][131] 	= partial_clause_prev[0][131] & x[50];
			partial_clause[0][132] 	= partial_clause_prev[0][132] & ~x[15] & ~x[44] & ~x[47] & ~x[59];
			partial_clause[0][133] 	= partial_clause_prev[0][133] & 1'b1;
			partial_clause[0][134] 	= partial_clause_prev[0][134] & 1'b1;
			partial_clause[0][135] 	= partial_clause_prev[0][135] & 1'b1;
			partial_clause[0][136] 	= partial_clause_prev[0][136] & ~x[14] & ~x[43];
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & 1'b1;
			partial_clause[0][139] 	= partial_clause_prev[0][139] & 1'b1;
			partial_clause[0][140] 	= partial_clause_prev[0][140] & 1'b1;
			partial_clause[0][141] 	= partial_clause_prev[0][141] & 1'b1;
			partial_clause[0][142] 	= partial_clause_prev[0][142] & 1'b1;
			partial_clause[0][143] 	= partial_clause_prev[0][143] & 1'b1;
			partial_clause[0][144] 	= partial_clause_prev[0][144] & 1'b1;
			partial_clause[0][145] 	= partial_clause_prev[0][145] & 1'b1;
			partial_clause[0][146] 	= partial_clause_prev[0][146] & x[50];
			partial_clause[0][147] 	= partial_clause_prev[0][147] & 1'b1;
			partial_clause[0][148] 	= partial_clause_prev[0][148] & 1'b1;
			partial_clause[0][149] 	= partial_clause_prev[0][149] & 1'b1;
			partial_clause[0][150] 	= partial_clause_prev[0][150] & 1'b1;
			partial_clause[0][151] 	= partial_clause_prev[0][151] & 1'b1;
			partial_clause[0][152] 	= partial_clause_prev[0][152] & 1'b1;
			partial_clause[0][153] 	= partial_clause_prev[0][153] & 1'b1;
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & 1'b1;
			partial_clause[0][156] 	= partial_clause_prev[0][156] & 1'b1;
			partial_clause[0][157] 	= partial_clause_prev[0][157] & 1'b1;
			partial_clause[0][158] 	= partial_clause_prev[0][158] & 1'b1;
			partial_clause[0][159] 	= partial_clause_prev[0][159] & 1'b1;
			partial_clause[0][160] 	= partial_clause_prev[0][160] & 1'b1;
			partial_clause[0][161] 	= partial_clause_prev[0][161] & 1'b1;
			partial_clause[0][162] 	= partial_clause_prev[0][162] & 1'b1;
			partial_clause[0][163] 	= partial_clause_prev[0][163] & 1'b1;
			partial_clause[0][164] 	= partial_clause_prev[0][164] & ~x[43];
			partial_clause[0][165] 	= partial_clause_prev[0][165] & 1'b1;
			partial_clause[0][166] 	= partial_clause_prev[0][166] & 1'b1;
			partial_clause[0][167] 	= partial_clause_prev[0][167] & 1'b1;
			partial_clause[0][168] 	= partial_clause_prev[0][168] & 1'b1;
			partial_clause[0][169] 	= partial_clause_prev[0][169] & x[50];
			partial_clause[0][170] 	= partial_clause_prev[0][170] & x[22];
			partial_clause[0][171] 	= partial_clause_prev[0][171] & 1'b1;
			partial_clause[0][172] 	= partial_clause_prev[0][172] & 1'b1;
			partial_clause[0][173] 	= partial_clause_prev[0][173] & 1'b1;
			partial_clause[0][174] 	= partial_clause_prev[0][174] & 1'b1;
			partial_clause[0][175] 	= partial_clause_prev[0][175] & 1'b1;
			partial_clause[0][176] 	= partial_clause_prev[0][176] & 1'b1;
			partial_clause[0][177] 	= partial_clause_prev[0][177] & 1'b1;
			partial_clause[0][178] 	= partial_clause_prev[0][178] & 1'b1;
			partial_clause[0][179] 	= partial_clause_prev[0][179] & ~x[19];
			partial_clause[0][180] 	= partial_clause_prev[0][180] & 1'b1;
			partial_clause[0][181] 	= partial_clause_prev[0][181] & 1'b1;
			partial_clause[0][182] 	= partial_clause_prev[0][182] & x[20] & x[22];
			partial_clause[0][183] 	= partial_clause_prev[0][183] & ~x[41] & ~x[43] & ~x[44];
			partial_clause[0][184] 	= partial_clause_prev[0][184] & 1'b1;
			partial_clause[0][185] 	= partial_clause_prev[0][185] & 1'b1;
			partial_clause[0][186] 	= partial_clause_prev[0][186] & 1'b1;
			partial_clause[0][187] 	= partial_clause_prev[0][187] & x[24];
			partial_clause[0][188] 	= partial_clause_prev[0][188] & 1'b1;
			partial_clause[0][189] 	= partial_clause_prev[0][189] & 1'b1;
			partial_clause[0][190] 	= partial_clause_prev[0][190] & 1'b1;
			partial_clause[0][191] 	= partial_clause_prev[0][191] & x[20] & x[22];
			partial_clause[0][192] 	= partial_clause_prev[0][192] & x[48] & x[50];
			partial_clause[0][193] 	= partial_clause_prev[0][193] & x[24];
			partial_clause[0][194] 	= partial_clause_prev[0][194] & 1'b1;
			partial_clause[0][195] 	= partial_clause_prev[0][195] & 1'b1;
			partial_clause[0][196] 	= partial_clause_prev[0][196] & 1'b1;
			partial_clause[0][197] 	= partial_clause_prev[0][197] & 1'b1;
			partial_clause[0][198] 	= partial_clause_prev[0][198] & 1'b1;
			partial_clause[0][199] 	= partial_clause_prev[0][199] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[54];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & x[22];
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & ~x[19];
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & x[50];
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & ~x[19] & x[50];
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & x[22];
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & 1'b1;
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & ~x[53];
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & x[49];
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & x[36];
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & 1'b1;
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & x[49];
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & x[49];
			partial_clause[1][99] 	= partial_clause_prev[1][99] & x[33];
			partial_clause[1][100] 	= partial_clause_prev[1][100] & 1'b1;
			partial_clause[1][101] 	= partial_clause_prev[1][101] & 1'b1;
			partial_clause[1][102] 	= partial_clause_prev[1][102] & 1'b1;
			partial_clause[1][103] 	= partial_clause_prev[1][103] & 1'b1;
			partial_clause[1][104] 	= partial_clause_prev[1][104] & x[18];
			partial_clause[1][105] 	= partial_clause_prev[1][105] & 1'b1;
			partial_clause[1][106] 	= partial_clause_prev[1][106] & 1'b1;
			partial_clause[1][107] 	= partial_clause_prev[1][107] & 1'b1;
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & 1'b1;
			partial_clause[1][110] 	= partial_clause_prev[1][110] & 1'b1;
			partial_clause[1][111] 	= partial_clause_prev[1][111] & 1'b1;
			partial_clause[1][112] 	= partial_clause_prev[1][112] & 1'b1;
			partial_clause[1][113] 	= partial_clause_prev[1][113] & 1'b1;
			partial_clause[1][114] 	= partial_clause_prev[1][114] & 1'b1;
			partial_clause[1][115] 	= partial_clause_prev[1][115] & ~x[50] & ~x[51];
			partial_clause[1][116] 	= partial_clause_prev[1][116] & 1'b1;
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & 1'b1;
			partial_clause[1][119] 	= partial_clause_prev[1][119] & 1'b1;
			partial_clause[1][120] 	= partial_clause_prev[1][120] & 1'b1;
			partial_clause[1][121] 	= partial_clause_prev[1][121] & 1'b1;
			partial_clause[1][122] 	= partial_clause_prev[1][122] & 1'b1;
			partial_clause[1][123] 	= partial_clause_prev[1][123] & 1'b1;
			partial_clause[1][124] 	= partial_clause_prev[1][124] & 1'b1;
			partial_clause[1][125] 	= partial_clause_prev[1][125] & x[53];
			partial_clause[1][126] 	= partial_clause_prev[1][126] & x[54];
			partial_clause[1][127] 	= partial_clause_prev[1][127] & 1'b1;
			partial_clause[1][128] 	= partial_clause_prev[1][128] & x[48];
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & 1'b1;
			partial_clause[1][131] 	= partial_clause_prev[1][131] & 1'b1;
			partial_clause[1][132] 	= partial_clause_prev[1][132] & x[46];
			partial_clause[1][133] 	= partial_clause_prev[1][133] & 1'b1;
			partial_clause[1][134] 	= partial_clause_prev[1][134] & 1'b1;
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & 1'b1;
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & 1'b1;
			partial_clause[1][139] 	= partial_clause_prev[1][139] & 1'b1;
			partial_clause[1][140] 	= partial_clause_prev[1][140] & 1'b1;
			partial_clause[1][141] 	= partial_clause_prev[1][141] & x[55];
			partial_clause[1][142] 	= partial_clause_prev[1][142] & 1'b1;
			partial_clause[1][143] 	= partial_clause_prev[1][143] & x[45];
			partial_clause[1][144] 	= partial_clause_prev[1][144] & 1'b1;
			partial_clause[1][145] 	= partial_clause_prev[1][145] & x[24];
			partial_clause[1][146] 	= partial_clause_prev[1][146] & 1'b1;
			partial_clause[1][147] 	= partial_clause_prev[1][147] & 1'b1;
			partial_clause[1][148] 	= partial_clause_prev[1][148] & x[46];
			partial_clause[1][149] 	= partial_clause_prev[1][149] & 1'b1;
			partial_clause[1][150] 	= partial_clause_prev[1][150] & 1'b1;
			partial_clause[1][151] 	= partial_clause_prev[1][151] & 1'b1;
			partial_clause[1][152] 	= partial_clause_prev[1][152] & 1'b1;
			partial_clause[1][153] 	= partial_clause_prev[1][153] & 1'b1;
			partial_clause[1][154] 	= partial_clause_prev[1][154] & 1'b1;
			partial_clause[1][155] 	= partial_clause_prev[1][155] & 1'b1;
			partial_clause[1][156] 	= partial_clause_prev[1][156] & 1'b1;
			partial_clause[1][157] 	= partial_clause_prev[1][157] & 1'b1;
			partial_clause[1][158] 	= partial_clause_prev[1][158] & 1'b1;
			partial_clause[1][159] 	= partial_clause_prev[1][159] & 1'b1;
			partial_clause[1][160] 	= partial_clause_prev[1][160] & 1'b1;
			partial_clause[1][161] 	= partial_clause_prev[1][161] & 1'b1;
			partial_clause[1][162] 	= partial_clause_prev[1][162] & 1'b1;
			partial_clause[1][163] 	= partial_clause_prev[1][163] & 1'b1;
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & 1'b1;
			partial_clause[1][166] 	= partial_clause_prev[1][166] & 1'b1;
			partial_clause[1][167] 	= partial_clause_prev[1][167] & 1'b1;
			partial_clause[1][168] 	= partial_clause_prev[1][168] & 1'b1;
			partial_clause[1][169] 	= partial_clause_prev[1][169] & x[54];
			partial_clause[1][170] 	= partial_clause_prev[1][170] & 1'b1;
			partial_clause[1][171] 	= partial_clause_prev[1][171] & x[19];
			partial_clause[1][172] 	= partial_clause_prev[1][172] & 1'b1;
			partial_clause[1][173] 	= partial_clause_prev[1][173] & 1'b1;
			partial_clause[1][174] 	= partial_clause_prev[1][174] & 1'b1;
			partial_clause[1][175] 	= partial_clause_prev[1][175] & 1'b1;
			partial_clause[1][176] 	= partial_clause_prev[1][176] & 1'b1;
			partial_clause[1][177] 	= partial_clause_prev[1][177] & 1'b1;
			partial_clause[1][178] 	= partial_clause_prev[1][178] & 1'b1;
			partial_clause[1][179] 	= partial_clause_prev[1][179] & 1'b1;
			partial_clause[1][180] 	= partial_clause_prev[1][180] & 1'b1;
			partial_clause[1][181] 	= partial_clause_prev[1][181] & 1'b1;
			partial_clause[1][182] 	= partial_clause_prev[1][182] & x[46];
			partial_clause[1][183] 	= partial_clause_prev[1][183] & 1'b1;
			partial_clause[1][184] 	= partial_clause_prev[1][184] & 1'b1;
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & 1'b1;
			partial_clause[1][187] 	= partial_clause_prev[1][187] & 1'b1;
			partial_clause[1][188] 	= partial_clause_prev[1][188] & 1'b1;
			partial_clause[1][189] 	= partial_clause_prev[1][189] & 1'b1;
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & 1'b1;
			partial_clause[1][192] 	= partial_clause_prev[1][192] & 1'b1;
			partial_clause[1][193] 	= partial_clause_prev[1][193] & 1'b1;
			partial_clause[1][194] 	= partial_clause_prev[1][194] & ~x[51];
			partial_clause[1][195] 	= partial_clause_prev[1][195] & 1'b1;
			partial_clause[1][196] 	= partial_clause_prev[1][196] & 1'b1;
			partial_clause[1][197] 	= partial_clause_prev[1][197] & 1'b1;
			partial_clause[1][198] 	= partial_clause_prev[1][198] & 1'b1;
			partial_clause[1][199] 	= partial_clause_prev[1][199] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & ~x[15] & ~x[17];
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & x[62];
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & ~x[31] & ~x[59];
			partial_clause[2][18] 	= partial_clause_prev[2][18] & ~x[15];
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & ~x[15];
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & ~x[16] & ~x[42];
			partial_clause[2][39] 	= partial_clause_prev[2][39] & ~x[14];
			partial_clause[2][40] 	= partial_clause_prev[2][40] & ~x[57];
			partial_clause[2][41] 	= partial_clause_prev[2][41] & ~x[1];
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & ~x[30] & ~x[56];
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & x[6];
			partial_clause[2][54] 	= partial_clause_prev[2][54] & x[47];
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & x[21];
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & ~x[31] & ~x[57];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & ~x[30];
			partial_clause[2][70] 	= partial_clause_prev[2][70] & ~x[17] & ~x[42];
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & x[33];
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & ~x[14] & ~x[15] & ~x[18];
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & x[19];
			partial_clause[2][84] 	= partial_clause_prev[2][84] & x[6];
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & ~x[43];
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & ~x[57];
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			partial_clause[2][100] 	= partial_clause_prev[2][100] & 1'b1;
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & ~x[45];
			partial_clause[2][103] 	= partial_clause_prev[2][103] & 1'b1;
			partial_clause[2][104] 	= partial_clause_prev[2][104] & 1'b1;
			partial_clause[2][105] 	= partial_clause_prev[2][105] & 1'b1;
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & 1'b1;
			partial_clause[2][108] 	= partial_clause_prev[2][108] & 1'b1;
			partial_clause[2][109] 	= partial_clause_prev[2][109] & 1'b1;
			partial_clause[2][110] 	= partial_clause_prev[2][110] & 1'b1;
			partial_clause[2][111] 	= partial_clause_prev[2][111] & 1'b1;
			partial_clause[2][112] 	= partial_clause_prev[2][112] & ~x[15];
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & ~x[15] & ~x[43];
			partial_clause[2][115] 	= partial_clause_prev[2][115] & 1'b1;
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & x[15];
			partial_clause[2][118] 	= partial_clause_prev[2][118] & ~x[59];
			partial_clause[2][119] 	= partial_clause_prev[2][119] & x[17];
			partial_clause[2][120] 	= partial_clause_prev[2][120] & 1'b1;
			partial_clause[2][121] 	= partial_clause_prev[2][121] & 1'b1;
			partial_clause[2][122] 	= partial_clause_prev[2][122] & x[43];
			partial_clause[2][123] 	= partial_clause_prev[2][123] & ~x[42];
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & 1'b1;
			partial_clause[2][126] 	= partial_clause_prev[2][126] & x[43];
			partial_clause[2][127] 	= partial_clause_prev[2][127] & 1'b1;
			partial_clause[2][128] 	= partial_clause_prev[2][128] & 1'b1;
			partial_clause[2][129] 	= partial_clause_prev[2][129] & 1'b1;
			partial_clause[2][130] 	= partial_clause_prev[2][130] & 1'b1;
			partial_clause[2][131] 	= partial_clause_prev[2][131] & ~x[15] & ~x[31];
			partial_clause[2][132] 	= partial_clause_prev[2][132] & x[45];
			partial_clause[2][133] 	= partial_clause_prev[2][133] & 1'b1;
			partial_clause[2][134] 	= partial_clause_prev[2][134] & 1'b1;
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & 1'b1;
			partial_clause[2][137] 	= partial_clause_prev[2][137] & 1'b1;
			partial_clause[2][138] 	= partial_clause_prev[2][138] & 1'b1;
			partial_clause[2][139] 	= partial_clause_prev[2][139] & 1'b1;
			partial_clause[2][140] 	= partial_clause_prev[2][140] & 1'b1;
			partial_clause[2][141] 	= partial_clause_prev[2][141] & x[19];
			partial_clause[2][142] 	= partial_clause_prev[2][142] & 1'b1;
			partial_clause[2][143] 	= partial_clause_prev[2][143] & 1'b1;
			partial_clause[2][144] 	= partial_clause_prev[2][144] & 1'b1;
			partial_clause[2][145] 	= partial_clause_prev[2][145] & 1'b1;
			partial_clause[2][146] 	= partial_clause_prev[2][146] & x[18];
			partial_clause[2][147] 	= partial_clause_prev[2][147] & 1'b1;
			partial_clause[2][148] 	= partial_clause_prev[2][148] & 1'b1;
			partial_clause[2][149] 	= partial_clause_prev[2][149] & 1'b1;
			partial_clause[2][150] 	= partial_clause_prev[2][150] & 1'b1;
			partial_clause[2][151] 	= partial_clause_prev[2][151] & 1'b1;
			partial_clause[2][152] 	= partial_clause_prev[2][152] & 1'b1;
			partial_clause[2][153] 	= partial_clause_prev[2][153] & 1'b1;
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & ~x[31];
			partial_clause[2][156] 	= partial_clause_prev[2][156] & 1'b1;
			partial_clause[2][157] 	= partial_clause_prev[2][157] & x[17];
			partial_clause[2][158] 	= partial_clause_prev[2][158] & 1'b1;
			partial_clause[2][159] 	= partial_clause_prev[2][159] & 1'b1;
			partial_clause[2][160] 	= partial_clause_prev[2][160] & 1'b1;
			partial_clause[2][161] 	= partial_clause_prev[2][161] & 1'b1;
			partial_clause[2][162] 	= partial_clause_prev[2][162] & 1'b1;
			partial_clause[2][163] 	= partial_clause_prev[2][163] & 1'b1;
			partial_clause[2][164] 	= partial_clause_prev[2][164] & x[46];
			partial_clause[2][165] 	= partial_clause_prev[2][165] & x[35];
			partial_clause[2][166] 	= partial_clause_prev[2][166] & 1'b1;
			partial_clause[2][167] 	= partial_clause_prev[2][167] & 1'b1;
			partial_clause[2][168] 	= partial_clause_prev[2][168] & 1'b1;
			partial_clause[2][169] 	= partial_clause_prev[2][169] & ~x[14];
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & 1'b1;
			partial_clause[2][173] 	= partial_clause_prev[2][173] & x[15];
			partial_clause[2][174] 	= partial_clause_prev[2][174] & x[16];
			partial_clause[2][175] 	= partial_clause_prev[2][175] & 1'b1;
			partial_clause[2][176] 	= partial_clause_prev[2][176] & 1'b1;
			partial_clause[2][177] 	= partial_clause_prev[2][177] & 1'b1;
			partial_clause[2][178] 	= partial_clause_prev[2][178] & ~x[59];
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & 1'b1;
			partial_clause[2][181] 	= partial_clause_prev[2][181] & ~x[60];
			partial_clause[2][182] 	= partial_clause_prev[2][182] & 1'b1;
			partial_clause[2][183] 	= partial_clause_prev[2][183] & 1'b1;
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & 1'b1;
			partial_clause[2][186] 	= partial_clause_prev[2][186] & 1'b1;
			partial_clause[2][187] 	= partial_clause_prev[2][187] & 1'b1;
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & 1'b1;
			partial_clause[2][190] 	= partial_clause_prev[2][190] & 1'b1;
			partial_clause[2][191] 	= partial_clause_prev[2][191] & 1'b1;
			partial_clause[2][192] 	= partial_clause_prev[2][192] & 1'b1;
			partial_clause[2][193] 	= partial_clause_prev[2][193] & 1'b1;
			partial_clause[2][194] 	= partial_clause_prev[2][194] & 1'b1;
			partial_clause[2][195] 	= partial_clause_prev[2][195] & 1'b1;
			partial_clause[2][196] 	= partial_clause_prev[2][196] & 1'b1;
			partial_clause[2][197] 	= partial_clause_prev[2][197] & 1'b1;
			partial_clause[2][198] 	= partial_clause_prev[2][198] & 1'b1;
			partial_clause[2][199] 	= partial_clause_prev[2][199] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & x[49];
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & x[48];
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & x[40];
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & x[55];
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & x[21];
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & 1'b1;
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & x[20];
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & ~x[47];
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & x[57];
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & x[20];
			partial_clause[3][96] 	= partial_clause_prev[3][96] & x[49];
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & ~x[47];
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			partial_clause[3][100] 	= partial_clause_prev[3][100] & 1'b1;
			partial_clause[3][101] 	= partial_clause_prev[3][101] & 1'b1;
			partial_clause[3][102] 	= partial_clause_prev[3][102] & 1'b1;
			partial_clause[3][103] 	= partial_clause_prev[3][103] & x[14];
			partial_clause[3][104] 	= partial_clause_prev[3][104] & x[3];
			partial_clause[3][105] 	= partial_clause_prev[3][105] & 1'b1;
			partial_clause[3][106] 	= partial_clause_prev[3][106] & ~x[26];
			partial_clause[3][107] 	= partial_clause_prev[3][107] & 1'b1;
			partial_clause[3][108] 	= partial_clause_prev[3][108] & 1'b1;
			partial_clause[3][109] 	= partial_clause_prev[3][109] & x[43];
			partial_clause[3][110] 	= partial_clause_prev[3][110] & 1'b1;
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & 1'b1;
			partial_clause[3][113] 	= partial_clause_prev[3][113] & 1'b1;
			partial_clause[3][114] 	= partial_clause_prev[3][114] & 1'b1;
			partial_clause[3][115] 	= partial_clause_prev[3][115] & x[17];
			partial_clause[3][116] 	= partial_clause_prev[3][116] & 1'b1;
			partial_clause[3][117] 	= partial_clause_prev[3][117] & x[4];
			partial_clause[3][118] 	= partial_clause_prev[3][118] & 1'b1;
			partial_clause[3][119] 	= partial_clause_prev[3][119] & 1'b1;
			partial_clause[3][120] 	= partial_clause_prev[3][120] & 1'b1;
			partial_clause[3][121] 	= partial_clause_prev[3][121] & 1'b1;
			partial_clause[3][122] 	= partial_clause_prev[3][122] & 1'b1;
			partial_clause[3][123] 	= partial_clause_prev[3][123] & 1'b1;
			partial_clause[3][124] 	= partial_clause_prev[3][124] & 1'b1;
			partial_clause[3][125] 	= partial_clause_prev[3][125] & 1'b1;
			partial_clause[3][126] 	= partial_clause_prev[3][126] & ~x[22];
			partial_clause[3][127] 	= partial_clause_prev[3][127] & 1'b1;
			partial_clause[3][128] 	= partial_clause_prev[3][128] & 1'b1;
			partial_clause[3][129] 	= partial_clause_prev[3][129] & 1'b1;
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & 1'b1;
			partial_clause[3][132] 	= partial_clause_prev[3][132] & 1'b1;
			partial_clause[3][133] 	= partial_clause_prev[3][133] & 1'b1;
			partial_clause[3][134] 	= partial_clause_prev[3][134] & 1'b1;
			partial_clause[3][135] 	= partial_clause_prev[3][135] & x[13];
			partial_clause[3][136] 	= partial_clause_prev[3][136] & 1'b1;
			partial_clause[3][137] 	= partial_clause_prev[3][137] & 1'b1;
			partial_clause[3][138] 	= partial_clause_prev[3][138] & 1'b1;
			partial_clause[3][139] 	= partial_clause_prev[3][139] & x[53];
			partial_clause[3][140] 	= partial_clause_prev[3][140] & x[15];
			partial_clause[3][141] 	= partial_clause_prev[3][141] & 1'b1;
			partial_clause[3][142] 	= partial_clause_prev[3][142] & 1'b1;
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & 1'b1;
			partial_clause[3][145] 	= partial_clause_prev[3][145] & 1'b1;
			partial_clause[3][146] 	= partial_clause_prev[3][146] & 1'b1;
			partial_clause[3][147] 	= partial_clause_prev[3][147] & ~x[21] & ~x[49];
			partial_clause[3][148] 	= partial_clause_prev[3][148] & x[1];
			partial_clause[3][149] 	= partial_clause_prev[3][149] & 1'b1;
			partial_clause[3][150] 	= partial_clause_prev[3][150] & 1'b1;
			partial_clause[3][151] 	= partial_clause_prev[3][151] & 1'b1;
			partial_clause[3][152] 	= partial_clause_prev[3][152] & ~x[55];
			partial_clause[3][153] 	= partial_clause_prev[3][153] & 1'b1;
			partial_clause[3][154] 	= partial_clause_prev[3][154] & 1'b1;
			partial_clause[3][155] 	= partial_clause_prev[3][155] & x[45];
			partial_clause[3][156] 	= partial_clause_prev[3][156] & 1'b1;
			partial_clause[3][157] 	= partial_clause_prev[3][157] & x[15];
			partial_clause[3][158] 	= partial_clause_prev[3][158] & 1'b1;
			partial_clause[3][159] 	= partial_clause_prev[3][159] & ~x[55];
			partial_clause[3][160] 	= partial_clause_prev[3][160] & 1'b1;
			partial_clause[3][161] 	= partial_clause_prev[3][161] & 1'b1;
			partial_clause[3][162] 	= partial_clause_prev[3][162] & 1'b1;
			partial_clause[3][163] 	= partial_clause_prev[3][163] & 1'b1;
			partial_clause[3][164] 	= partial_clause_prev[3][164] & x[47];
			partial_clause[3][165] 	= partial_clause_prev[3][165] & 1'b1;
			partial_clause[3][166] 	= partial_clause_prev[3][166] & 1'b1;
			partial_clause[3][167] 	= partial_clause_prev[3][167] & 1'b1;
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & 1'b1;
			partial_clause[3][170] 	= partial_clause_prev[3][170] & 1'b1;
			partial_clause[3][171] 	= partial_clause_prev[3][171] & 1'b1;
			partial_clause[3][172] 	= partial_clause_prev[3][172] & x[16];
			partial_clause[3][173] 	= partial_clause_prev[3][173] & 1'b1;
			partial_clause[3][174] 	= partial_clause_prev[3][174] & 1'b1;
			partial_clause[3][175] 	= partial_clause_prev[3][175] & 1'b1;
			partial_clause[3][176] 	= partial_clause_prev[3][176] & ~x[49];
			partial_clause[3][177] 	= partial_clause_prev[3][177] & 1'b1;
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & 1'b1;
			partial_clause[3][180] 	= partial_clause_prev[3][180] & 1'b1;
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & 1'b1;
			partial_clause[3][183] 	= partial_clause_prev[3][183] & 1'b1;
			partial_clause[3][184] 	= partial_clause_prev[3][184] & ~x[22];
			partial_clause[3][185] 	= partial_clause_prev[3][185] & 1'b1;
			partial_clause[3][186] 	= partial_clause_prev[3][186] & 1'b1;
			partial_clause[3][187] 	= partial_clause_prev[3][187] & 1'b1;
			partial_clause[3][188] 	= partial_clause_prev[3][188] & 1'b1;
			partial_clause[3][189] 	= partial_clause_prev[3][189] & x[49];
			partial_clause[3][190] 	= partial_clause_prev[3][190] & 1'b1;
			partial_clause[3][191] 	= partial_clause_prev[3][191] & ~x[19] & ~x[56];
			partial_clause[3][192] 	= partial_clause_prev[3][192] & 1'b1;
			partial_clause[3][193] 	= partial_clause_prev[3][193] & x[2];
			partial_clause[3][194] 	= partial_clause_prev[3][194] & 1'b1;
			partial_clause[3][195] 	= partial_clause_prev[3][195] & 1'b1;
			partial_clause[3][196] 	= partial_clause_prev[3][196] & 1'b1;
			partial_clause[3][197] 	= partial_clause_prev[3][197] & 1'b1;
			partial_clause[3][198] 	= partial_clause_prev[3][198] & 1'b1;
			partial_clause[3][199] 	= partial_clause_prev[3][199] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & x[41];
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & x[38];
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & x[18] & x[25];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & x[53];
			partial_clause[4][16] 	= partial_clause_prev[4][16] & x[6];
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & x[45];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & 1'b1;
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & x[17];
			partial_clause[4][35] 	= partial_clause_prev[4][35] & x[24];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & x[25];
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & 1'b1;
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & x[17] & x[54] & x[55];
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & x[52];
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & x[43];
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & x[18];
			partial_clause[4][80] 	= partial_clause_prev[4][80] & x[45];
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & x[45] & x[52];
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & x[43];
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & x[13];
			partial_clause[4][97] 	= partial_clause_prev[4][97] & x[15] & x[55];
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & x[17];
			partial_clause[4][100] 	= partial_clause_prev[4][100] & 1'b1;
			partial_clause[4][101] 	= partial_clause_prev[4][101] & 1'b1;
			partial_clause[4][102] 	= partial_clause_prev[4][102] & 1'b1;
			partial_clause[4][103] 	= partial_clause_prev[4][103] & 1'b1;
			partial_clause[4][104] 	= partial_clause_prev[4][104] & 1'b1;
			partial_clause[4][105] 	= partial_clause_prev[4][105] & 1'b1;
			partial_clause[4][106] 	= partial_clause_prev[4][106] & 1'b1;
			partial_clause[4][107] 	= partial_clause_prev[4][107] & 1'b1;
			partial_clause[4][108] 	= partial_clause_prev[4][108] & ~x[18];
			partial_clause[4][109] 	= partial_clause_prev[4][109] & 1'b1;
			partial_clause[4][110] 	= partial_clause_prev[4][110] & ~x[14];
			partial_clause[4][111] 	= partial_clause_prev[4][111] & 1'b1;
			partial_clause[4][112] 	= partial_clause_prev[4][112] & 1'b1;
			partial_clause[4][113] 	= partial_clause_prev[4][113] & 1'b1;
			partial_clause[4][114] 	= partial_clause_prev[4][114] & 1'b1;
			partial_clause[4][115] 	= partial_clause_prev[4][115] & 1'b1;
			partial_clause[4][116] 	= partial_clause_prev[4][116] & 1'b1;
			partial_clause[4][117] 	= partial_clause_prev[4][117] & ~x[19];
			partial_clause[4][118] 	= partial_clause_prev[4][118] & 1'b1;
			partial_clause[4][119] 	= partial_clause_prev[4][119] & 1'b1;
			partial_clause[4][120] 	= partial_clause_prev[4][120] & x[49] & ~x[53];
			partial_clause[4][121] 	= partial_clause_prev[4][121] & ~x[14] & ~x[56];
			partial_clause[4][122] 	= partial_clause_prev[4][122] & 1'b1;
			partial_clause[4][123] 	= partial_clause_prev[4][123] & 1'b1;
			partial_clause[4][124] 	= partial_clause_prev[4][124] & 1'b1;
			partial_clause[4][125] 	= partial_clause_prev[4][125] & 1'b1;
			partial_clause[4][126] 	= partial_clause_prev[4][126] & 1'b1;
			partial_clause[4][127] 	= partial_clause_prev[4][127] & ~x[51];
			partial_clause[4][128] 	= partial_clause_prev[4][128] & 1'b1;
			partial_clause[4][129] 	= partial_clause_prev[4][129] & 1'b1;
			partial_clause[4][130] 	= partial_clause_prev[4][130] & 1'b1;
			partial_clause[4][131] 	= partial_clause_prev[4][131] & 1'b1;
			partial_clause[4][132] 	= partial_clause_prev[4][132] & 1'b1;
			partial_clause[4][133] 	= partial_clause_prev[4][133] & 1'b1;
			partial_clause[4][134] 	= partial_clause_prev[4][134] & 1'b1;
			partial_clause[4][135] 	= partial_clause_prev[4][135] & ~x[20] & ~x[47];
			partial_clause[4][136] 	= partial_clause_prev[4][136] & 1'b1;
			partial_clause[4][137] 	= partial_clause_prev[4][137] & ~x[1] & ~x[17] & ~x[18];
			partial_clause[4][138] 	= partial_clause_prev[4][138] & ~x[14];
			partial_clause[4][139] 	= partial_clause_prev[4][139] & 1'b1;
			partial_clause[4][140] 	= partial_clause_prev[4][140] & ~x[43];
			partial_clause[4][141] 	= partial_clause_prev[4][141] & 1'b1;
			partial_clause[4][142] 	= partial_clause_prev[4][142] & 1'b1;
			partial_clause[4][143] 	= partial_clause_prev[4][143] & 1'b1;
			partial_clause[4][144] 	= partial_clause_prev[4][144] & ~x[58];
			partial_clause[4][145] 	= partial_clause_prev[4][145] & 1'b1;
			partial_clause[4][146] 	= partial_clause_prev[4][146] & 1'b1;
			partial_clause[4][147] 	= partial_clause_prev[4][147] & 1'b1;
			partial_clause[4][148] 	= partial_clause_prev[4][148] & 1'b1;
			partial_clause[4][149] 	= partial_clause_prev[4][149] & 1'b1;
			partial_clause[4][150] 	= partial_clause_prev[4][150] & ~x[46];
			partial_clause[4][151] 	= partial_clause_prev[4][151] & 1'b1;
			partial_clause[4][152] 	= partial_clause_prev[4][152] & 1'b1;
			partial_clause[4][153] 	= partial_clause_prev[4][153] & 1'b1;
			partial_clause[4][154] 	= partial_clause_prev[4][154] & 1'b1;
			partial_clause[4][155] 	= partial_clause_prev[4][155] & 1'b1;
			partial_clause[4][156] 	= partial_clause_prev[4][156] & ~x[25] & ~x[27];
			partial_clause[4][157] 	= partial_clause_prev[4][157] & 1'b1;
			partial_clause[4][158] 	= partial_clause_prev[4][158] & 1'b1;
			partial_clause[4][159] 	= partial_clause_prev[4][159] & ~x[44];
			partial_clause[4][160] 	= partial_clause_prev[4][160] & 1'b1;
			partial_clause[4][161] 	= partial_clause_prev[4][161] & ~x[19];
			partial_clause[4][162] 	= partial_clause_prev[4][162] & 1'b1;
			partial_clause[4][163] 	= partial_clause_prev[4][163] & 1'b1;
			partial_clause[4][164] 	= partial_clause_prev[4][164] & 1'b1;
			partial_clause[4][165] 	= partial_clause_prev[4][165] & 1'b1;
			partial_clause[4][166] 	= partial_clause_prev[4][166] & 1'b1;
			partial_clause[4][167] 	= partial_clause_prev[4][167] & 1'b1;
			partial_clause[4][168] 	= partial_clause_prev[4][168] & 1'b1;
			partial_clause[4][169] 	= partial_clause_prev[4][169] & 1'b1;
			partial_clause[4][170] 	= partial_clause_prev[4][170] & 1'b1;
			partial_clause[4][171] 	= partial_clause_prev[4][171] & 1'b1;
			partial_clause[4][172] 	= partial_clause_prev[4][172] & 1'b1;
			partial_clause[4][173] 	= partial_clause_prev[4][173] & 1'b1;
			partial_clause[4][174] 	= partial_clause_prev[4][174] & 1'b1;
			partial_clause[4][175] 	= partial_clause_prev[4][175] & 1'b1;
			partial_clause[4][176] 	= partial_clause_prev[4][176] & 1'b1;
			partial_clause[4][177] 	= partial_clause_prev[4][177] & 1'b1;
			partial_clause[4][178] 	= partial_clause_prev[4][178] & 1'b1;
			partial_clause[4][179] 	= partial_clause_prev[4][179] & 1'b1;
			partial_clause[4][180] 	= partial_clause_prev[4][180] & ~x[53];
			partial_clause[4][181] 	= partial_clause_prev[4][181] & 1'b1;
			partial_clause[4][182] 	= partial_clause_prev[4][182] & 1'b1;
			partial_clause[4][183] 	= partial_clause_prev[4][183] & 1'b1;
			partial_clause[4][184] 	= partial_clause_prev[4][184] & 1'b1;
			partial_clause[4][185] 	= partial_clause_prev[4][185] & 1'b1;
			partial_clause[4][186] 	= partial_clause_prev[4][186] & ~x[16];
			partial_clause[4][187] 	= partial_clause_prev[4][187] & 1'b1;
			partial_clause[4][188] 	= partial_clause_prev[4][188] & 1'b1;
			partial_clause[4][189] 	= partial_clause_prev[4][189] & ~x[25] & ~x[55];
			partial_clause[4][190] 	= partial_clause_prev[4][190] & 1'b1;
			partial_clause[4][191] 	= partial_clause_prev[4][191] & 1'b1;
			partial_clause[4][192] 	= partial_clause_prev[4][192] & 1'b1;
			partial_clause[4][193] 	= partial_clause_prev[4][193] & 1'b1;
			partial_clause[4][194] 	= partial_clause_prev[4][194] & ~x[14];
			partial_clause[4][195] 	= partial_clause_prev[4][195] & 1'b1;
			partial_clause[4][196] 	= partial_clause_prev[4][196] & 1'b1;
			partial_clause[4][197] 	= partial_clause_prev[4][197] & 1'b1;
			partial_clause[4][198] 	= partial_clause_prev[4][198] & 1'b1;
			partial_clause[4][199] 	= partial_clause_prev[4][199] & ~x[6] & ~x[41] & ~x[43];
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & ~x[52];
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & ~x[0] & ~x[4];
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & x[19];
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & ~x[56];
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & x[18] & ~x[55];
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & ~x[26];
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & ~x[43];
			partial_clause[5][69] 	= partial_clause_prev[5][69] & ~x[1];
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & ~x[13] & ~x[43];
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & ~x[27] & ~x[57];
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			partial_clause[5][100] 	= partial_clause_prev[5][100] & 1'b1;
			partial_clause[5][101] 	= partial_clause_prev[5][101] & 1'b1;
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & 1'b1;
			partial_clause[5][104] 	= partial_clause_prev[5][104] & 1'b1;
			partial_clause[5][105] 	= partial_clause_prev[5][105] & 1'b1;
			partial_clause[5][106] 	= partial_clause_prev[5][106] & 1'b1;
			partial_clause[5][107] 	= partial_clause_prev[5][107] & 1'b1;
			partial_clause[5][108] 	= partial_clause_prev[5][108] & x[61];
			partial_clause[5][109] 	= partial_clause_prev[5][109] & 1'b1;
			partial_clause[5][110] 	= partial_clause_prev[5][110] & 1'b1;
			partial_clause[5][111] 	= partial_clause_prev[5][111] & 1'b1;
			partial_clause[5][112] 	= partial_clause_prev[5][112] & 1'b1;
			partial_clause[5][113] 	= partial_clause_prev[5][113] & 1'b1;
			partial_clause[5][114] 	= partial_clause_prev[5][114] & x[4];
			partial_clause[5][115] 	= partial_clause_prev[5][115] & 1'b1;
			partial_clause[5][116] 	= partial_clause_prev[5][116] & 1'b1;
			partial_clause[5][117] 	= partial_clause_prev[5][117] & 1'b1;
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & 1'b1;
			partial_clause[5][120] 	= partial_clause_prev[5][120] & 1'b1;
			partial_clause[5][121] 	= partial_clause_prev[5][121] & 1'b1;
			partial_clause[5][122] 	= partial_clause_prev[5][122] & x[51];
			partial_clause[5][123] 	= partial_clause_prev[5][123] & 1'b1;
			partial_clause[5][124] 	= partial_clause_prev[5][124] & 1'b1;
			partial_clause[5][125] 	= partial_clause_prev[5][125] & ~x[0];
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & x[22];
			partial_clause[5][128] 	= partial_clause_prev[5][128] & 1'b1;
			partial_clause[5][129] 	= partial_clause_prev[5][129] & x[25];
			partial_clause[5][130] 	= partial_clause_prev[5][130] & 1'b1;
			partial_clause[5][131] 	= partial_clause_prev[5][131] & x[51];
			partial_clause[5][132] 	= partial_clause_prev[5][132] & 1'b1;
			partial_clause[5][133] 	= partial_clause_prev[5][133] & 1'b1;
			partial_clause[5][134] 	= partial_clause_prev[5][134] & 1'b1;
			partial_clause[5][135] 	= partial_clause_prev[5][135] & 1'b1;
			partial_clause[5][136] 	= partial_clause_prev[5][136] & 1'b1;
			partial_clause[5][137] 	= partial_clause_prev[5][137] & 1'b1;
			partial_clause[5][138] 	= partial_clause_prev[5][138] & 1'b1;
			partial_clause[5][139] 	= partial_clause_prev[5][139] & 1'b1;
			partial_clause[5][140] 	= partial_clause_prev[5][140] & x[0];
			partial_clause[5][141] 	= partial_clause_prev[5][141] & 1'b1;
			partial_clause[5][142] 	= partial_clause_prev[5][142] & 1'b1;
			partial_clause[5][143] 	= partial_clause_prev[5][143] & 1'b1;
			partial_clause[5][144] 	= partial_clause_prev[5][144] & x[51];
			partial_clause[5][145] 	= partial_clause_prev[5][145] & x[2];
			partial_clause[5][146] 	= partial_clause_prev[5][146] & 1'b1;
			partial_clause[5][147] 	= partial_clause_prev[5][147] & 1'b1;
			partial_clause[5][148] 	= partial_clause_prev[5][148] & 1'b1;
			partial_clause[5][149] 	= partial_clause_prev[5][149] & 1'b1;
			partial_clause[5][150] 	= partial_clause_prev[5][150] & 1'b1;
			partial_clause[5][151] 	= partial_clause_prev[5][151] & 1'b1;
			partial_clause[5][152] 	= partial_clause_prev[5][152] & 1'b1;
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & x[43];
			partial_clause[5][155] 	= partial_clause_prev[5][155] & 1'b1;
			partial_clause[5][156] 	= partial_clause_prev[5][156] & 1'b1;
			partial_clause[5][157] 	= partial_clause_prev[5][157] & 1'b1;
			partial_clause[5][158] 	= partial_clause_prev[5][158] & x[23];
			partial_clause[5][159] 	= partial_clause_prev[5][159] & 1'b1;
			partial_clause[5][160] 	= partial_clause_prev[5][160] & 1'b1;
			partial_clause[5][161] 	= partial_clause_prev[5][161] & ~x[18];
			partial_clause[5][162] 	= partial_clause_prev[5][162] & 1'b1;
			partial_clause[5][163] 	= partial_clause_prev[5][163] & 1'b1;
			partial_clause[5][164] 	= partial_clause_prev[5][164] & 1'b1;
			partial_clause[5][165] 	= partial_clause_prev[5][165] & 1'b1;
			partial_clause[5][166] 	= partial_clause_prev[5][166] & x[30];
			partial_clause[5][167] 	= partial_clause_prev[5][167] & 1'b1;
			partial_clause[5][168] 	= partial_clause_prev[5][168] & 1'b1;
			partial_clause[5][169] 	= partial_clause_prev[5][169] & 1'b1;
			partial_clause[5][170] 	= partial_clause_prev[5][170] & x[3];
			partial_clause[5][171] 	= partial_clause_prev[5][171] & 1'b1;
			partial_clause[5][172] 	= partial_clause_prev[5][172] & x[1];
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & 1'b1;
			partial_clause[5][175] 	= partial_clause_prev[5][175] & 1'b1;
			partial_clause[5][176] 	= partial_clause_prev[5][176] & x[42];
			partial_clause[5][177] 	= partial_clause_prev[5][177] & x[24];
			partial_clause[5][178] 	= partial_clause_prev[5][178] & 1'b1;
			partial_clause[5][179] 	= partial_clause_prev[5][179] & 1'b1;
			partial_clause[5][180] 	= partial_clause_prev[5][180] & x[51];
			partial_clause[5][181] 	= partial_clause_prev[5][181] & 1'b1;
			partial_clause[5][182] 	= partial_clause_prev[5][182] & x[25];
			partial_clause[5][183] 	= partial_clause_prev[5][183] & 1'b1;
			partial_clause[5][184] 	= partial_clause_prev[5][184] & x[29] & x[44];
			partial_clause[5][185] 	= partial_clause_prev[5][185] & 1'b1;
			partial_clause[5][186] 	= partial_clause_prev[5][186] & ~x[0];
			partial_clause[5][187] 	= partial_clause_prev[5][187] & 1'b1;
			partial_clause[5][188] 	= partial_clause_prev[5][188] & 1'b1;
			partial_clause[5][189] 	= partial_clause_prev[5][189] & 1'b1;
			partial_clause[5][190] 	= partial_clause_prev[5][190] & 1'b1;
			partial_clause[5][191] 	= partial_clause_prev[5][191] & 1'b1;
			partial_clause[5][192] 	= partial_clause_prev[5][192] & 1'b1;
			partial_clause[5][193] 	= partial_clause_prev[5][193] & x[50];
			partial_clause[5][194] 	= partial_clause_prev[5][194] & 1'b1;
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & 1'b1;
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & 1'b1;
			partial_clause[5][199] 	= partial_clause_prev[5][199] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & x[17];
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & x[30];
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & x[46];
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & x[19];
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & x[20] & x[47];
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & x[18];
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & x[61];
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & x[46];
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & x[30];
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & x[3] & x[31];
			partial_clause[6][76] 	= partial_clause_prev[6][76] & x[46];
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & ~x[54];
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & x[3];
			partial_clause[6][99] 	= partial_clause_prev[6][99] & x[42];
			partial_clause[6][100] 	= partial_clause_prev[6][100] & 1'b1;
			partial_clause[6][101] 	= partial_clause_prev[6][101] & 1'b1;
			partial_clause[6][102] 	= partial_clause_prev[6][102] & 1'b1;
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & 1'b1;
			partial_clause[6][105] 	= partial_clause_prev[6][105] & 1'b1;
			partial_clause[6][106] 	= partial_clause_prev[6][106] & ~x[2];
			partial_clause[6][107] 	= partial_clause_prev[6][107] & 1'b1;
			partial_clause[6][108] 	= partial_clause_prev[6][108] & ~x[44];
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & 1'b1;
			partial_clause[6][111] 	= partial_clause_prev[6][111] & 1'b1;
			partial_clause[6][112] 	= partial_clause_prev[6][112] & 1'b1;
			partial_clause[6][113] 	= partial_clause_prev[6][113] & ~x[58];
			partial_clause[6][114] 	= partial_clause_prev[6][114] & 1'b1;
			partial_clause[6][115] 	= partial_clause_prev[6][115] & 1'b1;
			partial_clause[6][116] 	= partial_clause_prev[6][116] & 1'b1;
			partial_clause[6][117] 	= partial_clause_prev[6][117] & 1'b1;
			partial_clause[6][118] 	= partial_clause_prev[6][118] & 1'b1;
			partial_clause[6][119] 	= partial_clause_prev[6][119] & 1'b1;
			partial_clause[6][120] 	= partial_clause_prev[6][120] & 1'b1;
			partial_clause[6][121] 	= partial_clause_prev[6][121] & ~x[15];
			partial_clause[6][122] 	= partial_clause_prev[6][122] & 1'b1;
			partial_clause[6][123] 	= partial_clause_prev[6][123] & 1'b1;
			partial_clause[6][124] 	= partial_clause_prev[6][124] & 1'b1;
			partial_clause[6][125] 	= partial_clause_prev[6][125] & ~x[47];
			partial_clause[6][126] 	= partial_clause_prev[6][126] & 1'b1;
			partial_clause[6][127] 	= partial_clause_prev[6][127] & 1'b1;
			partial_clause[6][128] 	= partial_clause_prev[6][128] & 1'b1;
			partial_clause[6][129] 	= partial_clause_prev[6][129] & 1'b1;
			partial_clause[6][130] 	= partial_clause_prev[6][130] & 1'b1;
			partial_clause[6][131] 	= partial_clause_prev[6][131] & 1'b1;
			partial_clause[6][132] 	= partial_clause_prev[6][132] & 1'b1;
			partial_clause[6][133] 	= partial_clause_prev[6][133] & 1'b1;
			partial_clause[6][134] 	= partial_clause_prev[6][134] & 1'b1;
			partial_clause[6][135] 	= partial_clause_prev[6][135] & 1'b1;
			partial_clause[6][136] 	= partial_clause_prev[6][136] & 1'b1;
			partial_clause[6][137] 	= partial_clause_prev[6][137] & 1'b1;
			partial_clause[6][138] 	= partial_clause_prev[6][138] & 1'b1;
			partial_clause[6][139] 	= partial_clause_prev[6][139] & 1'b1;
			partial_clause[6][140] 	= partial_clause_prev[6][140] & 1'b1;
			partial_clause[6][141] 	= partial_clause_prev[6][141] & 1'b1;
			partial_clause[6][142] 	= partial_clause_prev[6][142] & 1'b1;
			partial_clause[6][143] 	= partial_clause_prev[6][143] & 1'b1;
			partial_clause[6][144] 	= partial_clause_prev[6][144] & 1'b1;
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & 1'b1;
			partial_clause[6][147] 	= partial_clause_prev[6][147] & 1'b1;
			partial_clause[6][148] 	= partial_clause_prev[6][148] & 1'b1;
			partial_clause[6][149] 	= partial_clause_prev[6][149] & 1'b1;
			partial_clause[6][150] 	= partial_clause_prev[6][150] & 1'b1;
			partial_clause[6][151] 	= partial_clause_prev[6][151] & 1'b1;
			partial_clause[6][152] 	= partial_clause_prev[6][152] & 1'b1;
			partial_clause[6][153] 	= partial_clause_prev[6][153] & ~x[20] & ~x[51];
			partial_clause[6][154] 	= partial_clause_prev[6][154] & ~x[0];
			partial_clause[6][155] 	= partial_clause_prev[6][155] & ~x[24];
			partial_clause[6][156] 	= partial_clause_prev[6][156] & 1'b1;
			partial_clause[6][157] 	= partial_clause_prev[6][157] & 1'b1;
			partial_clause[6][158] 	= partial_clause_prev[6][158] & 1'b1;
			partial_clause[6][159] 	= partial_clause_prev[6][159] & 1'b1;
			partial_clause[6][160] 	= partial_clause_prev[6][160] & ~x[43];
			partial_clause[6][161] 	= partial_clause_prev[6][161] & 1'b1;
			partial_clause[6][162] 	= partial_clause_prev[6][162] & 1'b1;
			partial_clause[6][163] 	= partial_clause_prev[6][163] & 1'b1;
			partial_clause[6][164] 	= partial_clause_prev[6][164] & 1'b1;
			partial_clause[6][165] 	= partial_clause_prev[6][165] & 1'b1;
			partial_clause[6][166] 	= partial_clause_prev[6][166] & 1'b1;
			partial_clause[6][167] 	= partial_clause_prev[6][167] & 1'b1;
			partial_clause[6][168] 	= partial_clause_prev[6][168] & 1'b1;
			partial_clause[6][169] 	= partial_clause_prev[6][169] & ~x[31];
			partial_clause[6][170] 	= partial_clause_prev[6][170] & 1'b1;
			partial_clause[6][171] 	= partial_clause_prev[6][171] & 1'b1;
			partial_clause[6][172] 	= partial_clause_prev[6][172] & 1'b1;
			partial_clause[6][173] 	= partial_clause_prev[6][173] & 1'b1;
			partial_clause[6][174] 	= partial_clause_prev[6][174] & 1'b1;
			partial_clause[6][175] 	= partial_clause_prev[6][175] & 1'b1;
			partial_clause[6][176] 	= partial_clause_prev[6][176] & ~x[30] & ~x[31];
			partial_clause[6][177] 	= partial_clause_prev[6][177] & 1'b1;
			partial_clause[6][178] 	= partial_clause_prev[6][178] & 1'b1;
			partial_clause[6][179] 	= partial_clause_prev[6][179] & 1'b1;
			partial_clause[6][180] 	= partial_clause_prev[6][180] & 1'b1;
			partial_clause[6][181] 	= partial_clause_prev[6][181] & 1'b1;
			partial_clause[6][182] 	= partial_clause_prev[6][182] & 1'b1;
			partial_clause[6][183] 	= partial_clause_prev[6][183] & ~x[3] & ~x[14];
			partial_clause[6][184] 	= partial_clause_prev[6][184] & 1'b1;
			partial_clause[6][185] 	= partial_clause_prev[6][185] & 1'b1;
			partial_clause[6][186] 	= partial_clause_prev[6][186] & 1'b1;
			partial_clause[6][187] 	= partial_clause_prev[6][187] & 1'b1;
			partial_clause[6][188] 	= partial_clause_prev[6][188] & 1'b1;
			partial_clause[6][189] 	= partial_clause_prev[6][189] & 1'b1;
			partial_clause[6][190] 	= partial_clause_prev[6][190] & 1'b1;
			partial_clause[6][191] 	= partial_clause_prev[6][191] & 1'b1;
			partial_clause[6][192] 	= partial_clause_prev[6][192] & 1'b1;
			partial_clause[6][193] 	= partial_clause_prev[6][193] & ~x[3];
			partial_clause[6][194] 	= partial_clause_prev[6][194] & 1'b1;
			partial_clause[6][195] 	= partial_clause_prev[6][195] & 1'b1;
			partial_clause[6][196] 	= partial_clause_prev[6][196] & 1'b1;
			partial_clause[6][197] 	= partial_clause_prev[6][197] & 1'b1;
			partial_clause[6][198] 	= partial_clause_prev[6][198] & 1'b1;
			partial_clause[6][199] 	= partial_clause_prev[6][199] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & x[9];
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & ~x[49];
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & ~x[22];
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & ~x[47];
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & ~x[49] & ~x[50];
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & ~x[23];
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & x[39];
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & x[53];
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & x[51];
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & ~x[47];
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & ~x[22];
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & x[5];
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & ~x[21] & ~x[49];
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & ~x[29];
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & ~x[30] & ~x[48];
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & ~x[22] & ~x[49];
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			partial_clause[7][100] 	= partial_clause_prev[7][100] & ~x[53];
			partial_clause[7][101] 	= partial_clause_prev[7][101] & x[21] & ~x[55];
			partial_clause[7][102] 	= partial_clause_prev[7][102] & 1'b1;
			partial_clause[7][103] 	= partial_clause_prev[7][103] & 1'b1;
			partial_clause[7][104] 	= partial_clause_prev[7][104] & x[47];
			partial_clause[7][105] 	= partial_clause_prev[7][105] & 1'b1;
			partial_clause[7][106] 	= partial_clause_prev[7][106] & 1'b1;
			partial_clause[7][107] 	= partial_clause_prev[7][107] & 1'b1;
			partial_clause[7][108] 	= partial_clause_prev[7][108] & 1'b1;
			partial_clause[7][109] 	= partial_clause_prev[7][109] & 1'b1;
			partial_clause[7][110] 	= partial_clause_prev[7][110] & 1'b1;
			partial_clause[7][111] 	= partial_clause_prev[7][111] & 1'b1;
			partial_clause[7][112] 	= partial_clause_prev[7][112] & 1'b1;
			partial_clause[7][113] 	= partial_clause_prev[7][113] & 1'b1;
			partial_clause[7][114] 	= partial_clause_prev[7][114] & 1'b1;
			partial_clause[7][115] 	= partial_clause_prev[7][115] & 1'b1;
			partial_clause[7][116] 	= partial_clause_prev[7][116] & 1'b1;
			partial_clause[7][117] 	= partial_clause_prev[7][117] & 1'b1;
			partial_clause[7][118] 	= partial_clause_prev[7][118] & 1'b1;
			partial_clause[7][119] 	= partial_clause_prev[7][119] & 1'b1;
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & 1'b1;
			partial_clause[7][123] 	= partial_clause_prev[7][123] & 1'b1;
			partial_clause[7][124] 	= partial_clause_prev[7][124] & x[45];
			partial_clause[7][125] 	= partial_clause_prev[7][125] & 1'b1;
			partial_clause[7][126] 	= partial_clause_prev[7][126] & 1'b1;
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & 1'b1;
			partial_clause[7][129] 	= partial_clause_prev[7][129] & x[22] & ~x[57];
			partial_clause[7][130] 	= partial_clause_prev[7][130] & 1'b1;
			partial_clause[7][131] 	= partial_clause_prev[7][131] & x[21];
			partial_clause[7][132] 	= partial_clause_prev[7][132] & 1'b1;
			partial_clause[7][133] 	= partial_clause_prev[7][133] & x[43];
			partial_clause[7][134] 	= partial_clause_prev[7][134] & 1'b1;
			partial_clause[7][135] 	= partial_clause_prev[7][135] & 1'b1;
			partial_clause[7][136] 	= partial_clause_prev[7][136] & 1'b1;
			partial_clause[7][137] 	= partial_clause_prev[7][137] & ~x[33];
			partial_clause[7][138] 	= partial_clause_prev[7][138] & 1'b1;
			partial_clause[7][139] 	= partial_clause_prev[7][139] & x[17];
			partial_clause[7][140] 	= partial_clause_prev[7][140] & x[17] & x[50];
			partial_clause[7][141] 	= partial_clause_prev[7][141] & ~x[0];
			partial_clause[7][142] 	= partial_clause_prev[7][142] & x[48];
			partial_clause[7][143] 	= partial_clause_prev[7][143] & 1'b1;
			partial_clause[7][144] 	= partial_clause_prev[7][144] & 1'b1;
			partial_clause[7][145] 	= partial_clause_prev[7][145] & x[43];
			partial_clause[7][146] 	= partial_clause_prev[7][146] & x[21] & ~x[27];
			partial_clause[7][147] 	= partial_clause_prev[7][147] & x[16];
			partial_clause[7][148] 	= partial_clause_prev[7][148] & 1'b1;
			partial_clause[7][149] 	= partial_clause_prev[7][149] & 1'b1;
			partial_clause[7][150] 	= partial_clause_prev[7][150] & x[18];
			partial_clause[7][151] 	= partial_clause_prev[7][151] & x[15];
			partial_clause[7][152] 	= partial_clause_prev[7][152] & 1'b1;
			partial_clause[7][153] 	= partial_clause_prev[7][153] & x[48];
			partial_clause[7][154] 	= partial_clause_prev[7][154] & x[19] & x[48];
			partial_clause[7][155] 	= partial_clause_prev[7][155] & x[19] & ~x[56];
			partial_clause[7][156] 	= partial_clause_prev[7][156] & 1'b1;
			partial_clause[7][157] 	= partial_clause_prev[7][157] & x[19];
			partial_clause[7][158] 	= partial_clause_prev[7][158] & 1'b1;
			partial_clause[7][159] 	= partial_clause_prev[7][159] & 1'b1;
			partial_clause[7][160] 	= partial_clause_prev[7][160] & 1'b1;
			partial_clause[7][161] 	= partial_clause_prev[7][161] & 1'b1;
			partial_clause[7][162] 	= partial_clause_prev[7][162] & 1'b1;
			partial_clause[7][163] 	= partial_clause_prev[7][163] & 1'b1;
			partial_clause[7][164] 	= partial_clause_prev[7][164] & 1'b1;
			partial_clause[7][165] 	= partial_clause_prev[7][165] & 1'b1;
			partial_clause[7][166] 	= partial_clause_prev[7][166] & ~x[28];
			partial_clause[7][167] 	= partial_clause_prev[7][167] & 1'b1;
			partial_clause[7][168] 	= partial_clause_prev[7][168] & 1'b1;
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & ~x[1];
			partial_clause[7][171] 	= partial_clause_prev[7][171] & x[20] & ~x[28];
			partial_clause[7][172] 	= partial_clause_prev[7][172] & x[21] & ~x[30];
			partial_clause[7][173] 	= partial_clause_prev[7][173] & 1'b1;
			partial_clause[7][174] 	= partial_clause_prev[7][174] & 1'b1;
			partial_clause[7][175] 	= partial_clause_prev[7][175] & 1'b1;
			partial_clause[7][176] 	= partial_clause_prev[7][176] & 1'b1;
			partial_clause[7][177] 	= partial_clause_prev[7][177] & 1'b1;
			partial_clause[7][178] 	= partial_clause_prev[7][178] & 1'b1;
			partial_clause[7][179] 	= partial_clause_prev[7][179] & x[21];
			partial_clause[7][180] 	= partial_clause_prev[7][180] & ~x[56];
			partial_clause[7][181] 	= partial_clause_prev[7][181] & x[20] & ~x[29];
			partial_clause[7][182] 	= partial_clause_prev[7][182] & 1'b1;
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & 1'b1;
			partial_clause[7][185] 	= partial_clause_prev[7][185] & 1'b1;
			partial_clause[7][186] 	= partial_clause_prev[7][186] & 1'b1;
			partial_clause[7][187] 	= partial_clause_prev[7][187] & x[17];
			partial_clause[7][188] 	= partial_clause_prev[7][188] & x[17] & x[45];
			partial_clause[7][189] 	= partial_clause_prev[7][189] & 1'b1;
			partial_clause[7][190] 	= partial_clause_prev[7][190] & ~x[29];
			partial_clause[7][191] 	= partial_clause_prev[7][191] & 1'b1;
			partial_clause[7][192] 	= partial_clause_prev[7][192] & 1'b1;
			partial_clause[7][193] 	= partial_clause_prev[7][193] & ~x[56];
			partial_clause[7][194] 	= partial_clause_prev[7][194] & 1'b1;
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & ~x[0];
			partial_clause[7][197] 	= partial_clause_prev[7][197] & x[16];
			partial_clause[7][198] 	= partial_clause_prev[7][198] & 1'b1;
			partial_clause[7][199] 	= partial_clause_prev[7][199] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & x[39];
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & ~x[16] & x[48];
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & ~x[63];
			partial_clause[8][12] 	= partial_clause_prev[8][12] & ~x[45];
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & x[22] & ~x[26] & ~x[55];
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & x[51];
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & x[50];
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & ~x[2];
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & ~x[17] & x[21];
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & x[36];
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & ~x[27];
			partial_clause[8][56] 	= partial_clause_prev[8][56] & x[49];
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & ~x[16] & x[49];
			partial_clause[8][69] 	= partial_clause_prev[8][69] & ~x[57];
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & ~x[18] & x[50];
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & ~x[15] & ~x[44];
			partial_clause[8][82] 	= partial_clause_prev[8][82] & ~x[12];
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & ~x[56];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			partial_clause[8][100] 	= partial_clause_prev[8][100] & 1'b1;
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & 1'b1;
			partial_clause[8][103] 	= partial_clause_prev[8][103] & x[56];
			partial_clause[8][104] 	= partial_clause_prev[8][104] & 1'b1;
			partial_clause[8][105] 	= partial_clause_prev[8][105] & 1'b1;
			partial_clause[8][106] 	= partial_clause_prev[8][106] & 1'b1;
			partial_clause[8][107] 	= partial_clause_prev[8][107] & ~x[19];
			partial_clause[8][108] 	= partial_clause_prev[8][108] & 1'b1;
			partial_clause[8][109] 	= partial_clause_prev[8][109] & 1'b1;
			partial_clause[8][110] 	= partial_clause_prev[8][110] & 1'b1;
			partial_clause[8][111] 	= partial_clause_prev[8][111] & 1'b1;
			partial_clause[8][112] 	= partial_clause_prev[8][112] & ~x[20] & ~x[47];
			partial_clause[8][113] 	= partial_clause_prev[8][113] & 1'b1;
			partial_clause[8][114] 	= partial_clause_prev[8][114] & 1'b1;
			partial_clause[8][115] 	= partial_clause_prev[8][115] & 1'b1;
			partial_clause[8][116] 	= partial_clause_prev[8][116] & 1'b1;
			partial_clause[8][117] 	= partial_clause_prev[8][117] & 1'b1;
			partial_clause[8][118] 	= partial_clause_prev[8][118] & 1'b1;
			partial_clause[8][119] 	= partial_clause_prev[8][119] & 1'b1;
			partial_clause[8][120] 	= partial_clause_prev[8][120] & x[42];
			partial_clause[8][121] 	= partial_clause_prev[8][121] & 1'b1;
			partial_clause[8][122] 	= partial_clause_prev[8][122] & 1'b1;
			partial_clause[8][123] 	= partial_clause_prev[8][123] & 1'b1;
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & 1'b1;
			partial_clause[8][126] 	= partial_clause_prev[8][126] & x[55];
			partial_clause[8][127] 	= partial_clause_prev[8][127] & 1'b1;
			partial_clause[8][128] 	= partial_clause_prev[8][128] & 1'b1;
			partial_clause[8][129] 	= partial_clause_prev[8][129] & 1'b1;
			partial_clause[8][130] 	= partial_clause_prev[8][130] & 1'b1;
			partial_clause[8][131] 	= partial_clause_prev[8][131] & 1'b1;
			partial_clause[8][132] 	= partial_clause_prev[8][132] & 1'b1;
			partial_clause[8][133] 	= partial_clause_prev[8][133] & 1'b1;
			partial_clause[8][134] 	= partial_clause_prev[8][134] & 1'b1;
			partial_clause[8][135] 	= partial_clause_prev[8][135] & 1'b1;
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & 1'b1;
			partial_clause[8][138] 	= partial_clause_prev[8][138] & 1'b1;
			partial_clause[8][139] 	= partial_clause_prev[8][139] & 1'b1;
			partial_clause[8][140] 	= partial_clause_prev[8][140] & 1'b1;
			partial_clause[8][141] 	= partial_clause_prev[8][141] & 1'b1;
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & 1'b1;
			partial_clause[8][144] 	= partial_clause_prev[8][144] & 1'b1;
			partial_clause[8][145] 	= partial_clause_prev[8][145] & 1'b1;
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & x[59];
			partial_clause[8][148] 	= partial_clause_prev[8][148] & 1'b1;
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & 1'b1;
			partial_clause[8][151] 	= partial_clause_prev[8][151] & 1'b1;
			partial_clause[8][152] 	= partial_clause_prev[8][152] & 1'b1;
			partial_clause[8][153] 	= partial_clause_prev[8][153] & ~x[19];
			partial_clause[8][154] 	= partial_clause_prev[8][154] & x[60];
			partial_clause[8][155] 	= partial_clause_prev[8][155] & 1'b1;
			partial_clause[8][156] 	= partial_clause_prev[8][156] & ~x[21] & ~x[48];
			partial_clause[8][157] 	= partial_clause_prev[8][157] & 1'b1;
			partial_clause[8][158] 	= partial_clause_prev[8][158] & 1'b1;
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & 1'b1;
			partial_clause[8][161] 	= partial_clause_prev[8][161] & 1'b1;
			partial_clause[8][162] 	= partial_clause_prev[8][162] & x[44];
			partial_clause[8][163] 	= partial_clause_prev[8][163] & 1'b1;
			partial_clause[8][164] 	= partial_clause_prev[8][164] & ~x[18];
			partial_clause[8][165] 	= partial_clause_prev[8][165] & 1'b1;
			partial_clause[8][166] 	= partial_clause_prev[8][166] & 1'b1;
			partial_clause[8][167] 	= partial_clause_prev[8][167] & 1'b1;
			partial_clause[8][168] 	= partial_clause_prev[8][168] & ~x[49];
			partial_clause[8][169] 	= partial_clause_prev[8][169] & 1'b1;
			partial_clause[8][170] 	= partial_clause_prev[8][170] & 1'b1;
			partial_clause[8][171] 	= partial_clause_prev[8][171] & 1'b1;
			partial_clause[8][172] 	= partial_clause_prev[8][172] & x[41];
			partial_clause[8][173] 	= partial_clause_prev[8][173] & 1'b1;
			partial_clause[8][174] 	= partial_clause_prev[8][174] & 1'b1;
			partial_clause[8][175] 	= partial_clause_prev[8][175] & 1'b1;
			partial_clause[8][176] 	= partial_clause_prev[8][176] & 1'b1;
			partial_clause[8][177] 	= partial_clause_prev[8][177] & 1'b1;
			partial_clause[8][178] 	= partial_clause_prev[8][178] & 1'b1;
			partial_clause[8][179] 	= partial_clause_prev[8][179] & 1'b1;
			partial_clause[8][180] 	= partial_clause_prev[8][180] & 1'b1;
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & 1'b1;
			partial_clause[8][183] 	= partial_clause_prev[8][183] & ~x[21] & ~x[36] & ~x[48];
			partial_clause[8][184] 	= partial_clause_prev[8][184] & 1'b1;
			partial_clause[8][185] 	= partial_clause_prev[8][185] & 1'b1;
			partial_clause[8][186] 	= partial_clause_prev[8][186] & 1'b1;
			partial_clause[8][187] 	= partial_clause_prev[8][187] & 1'b1;
			partial_clause[8][188] 	= partial_clause_prev[8][188] & ~x[24] & ~x[52];
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & 1'b1;
			partial_clause[8][191] 	= partial_clause_prev[8][191] & 1'b1;
			partial_clause[8][192] 	= partial_clause_prev[8][192] & ~x[19] & ~x[53];
			partial_clause[8][193] 	= partial_clause_prev[8][193] & ~x[49] & ~x[50];
			partial_clause[8][194] 	= partial_clause_prev[8][194] & 1'b1;
			partial_clause[8][195] 	= partial_clause_prev[8][195] & 1'b1;
			partial_clause[8][196] 	= partial_clause_prev[8][196] & x[42];
			partial_clause[8][197] 	= partial_clause_prev[8][197] & 1'b1;
			partial_clause[8][198] 	= partial_clause_prev[8][198] & 1'b1;
			partial_clause[8][199] 	= partial_clause_prev[8][199] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & x[25];
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & x[25];
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & 1'b1;
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & x[13];
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & x[39];
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & x[21];
			partial_clause[9][69] 	= partial_clause_prev[9][69] & x[12];
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & x[47];
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & x[11];
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & ~x[19];
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & x[46] & ~x[56];
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & x[34];
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & x[16] & x[25];
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
			partial_clause[9][100] 	= partial_clause_prev[9][100] & ~x[24] & ~x[40];
			partial_clause[9][101] 	= partial_clause_prev[9][101] & 1'b1;
			partial_clause[9][102] 	= partial_clause_prev[9][102] & 1'b1;
			partial_clause[9][103] 	= partial_clause_prev[9][103] & 1'b1;
			partial_clause[9][104] 	= partial_clause_prev[9][104] & 1'b1;
			partial_clause[9][105] 	= partial_clause_prev[9][105] & 1'b1;
			partial_clause[9][106] 	= partial_clause_prev[9][106] & 1'b1;
			partial_clause[9][107] 	= partial_clause_prev[9][107] & 1'b1;
			partial_clause[9][108] 	= partial_clause_prev[9][108] & 1'b1;
			partial_clause[9][109] 	= partial_clause_prev[9][109] & 1'b1;
			partial_clause[9][110] 	= partial_clause_prev[9][110] & 1'b1;
			partial_clause[9][111] 	= partial_clause_prev[9][111] & ~x[11] & ~x[15] & ~x[42];
			partial_clause[9][112] 	= partial_clause_prev[9][112] & 1'b1;
			partial_clause[9][113] 	= partial_clause_prev[9][113] & 1'b1;
			partial_clause[9][114] 	= partial_clause_prev[9][114] & ~x[25];
			partial_clause[9][115] 	= partial_clause_prev[9][115] & 1'b1;
			partial_clause[9][116] 	= partial_clause_prev[9][116] & 1'b1;
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & 1'b1;
			partial_clause[9][119] 	= partial_clause_prev[9][119] & 1'b1;
			partial_clause[9][120] 	= partial_clause_prev[9][120] & 1'b1;
			partial_clause[9][121] 	= partial_clause_prev[9][121] & 1'b1;
			partial_clause[9][122] 	= partial_clause_prev[9][122] & 1'b1;
			partial_clause[9][123] 	= partial_clause_prev[9][123] & 1'b1;
			partial_clause[9][124] 	= partial_clause_prev[9][124] & 1'b1;
			partial_clause[9][125] 	= partial_clause_prev[9][125] & 1'b1;
			partial_clause[9][126] 	= partial_clause_prev[9][126] & 1'b1;
			partial_clause[9][127] 	= partial_clause_prev[9][127] & 1'b1;
			partial_clause[9][128] 	= partial_clause_prev[9][128] & 1'b1;
			partial_clause[9][129] 	= partial_clause_prev[9][129] & ~x[21] & ~x[49];
			partial_clause[9][130] 	= partial_clause_prev[9][130] & 1'b1;
			partial_clause[9][131] 	= partial_clause_prev[9][131] & 1'b1;
			partial_clause[9][132] 	= partial_clause_prev[9][132] & 1'b1;
			partial_clause[9][133] 	= partial_clause_prev[9][133] & 1'b1;
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & 1'b1;
			partial_clause[9][138] 	= partial_clause_prev[9][138] & 1'b1;
			partial_clause[9][139] 	= partial_clause_prev[9][139] & 1'b1;
			partial_clause[9][140] 	= partial_clause_prev[9][140] & 1'b1;
			partial_clause[9][141] 	= partial_clause_prev[9][141] & 1'b1;
			partial_clause[9][142] 	= partial_clause_prev[9][142] & 1'b1;
			partial_clause[9][143] 	= partial_clause_prev[9][143] & 1'b1;
			partial_clause[9][144] 	= partial_clause_prev[9][144] & 1'b1;
			partial_clause[9][145] 	= partial_clause_prev[9][145] & 1'b1;
			partial_clause[9][146] 	= partial_clause_prev[9][146] & 1'b1;
			partial_clause[9][147] 	= partial_clause_prev[9][147] & ~x[13];
			partial_clause[9][148] 	= partial_clause_prev[9][148] & ~x[18] & ~x[20] & ~x[45];
			partial_clause[9][149] 	= partial_clause_prev[9][149] & ~x[18] & ~x[41] & ~x[42] & ~x[44];
			partial_clause[9][150] 	= partial_clause_prev[9][150] & 1'b1;
			partial_clause[9][151] 	= partial_clause_prev[9][151] & x[49];
			partial_clause[9][152] 	= partial_clause_prev[9][152] & 1'b1;
			partial_clause[9][153] 	= partial_clause_prev[9][153] & 1'b1;
			partial_clause[9][154] 	= partial_clause_prev[9][154] & ~x[15] & ~x[16] & ~x[41];
			partial_clause[9][155] 	= partial_clause_prev[9][155] & 1'b1;
			partial_clause[9][156] 	= partial_clause_prev[9][156] & 1'b1;
			partial_clause[9][157] 	= partial_clause_prev[9][157] & ~x[1];
			partial_clause[9][158] 	= partial_clause_prev[9][158] & ~x[16] & ~x[41] & ~x[43];
			partial_clause[9][159] 	= partial_clause_prev[9][159] & 1'b1;
			partial_clause[9][160] 	= partial_clause_prev[9][160] & 1'b1;
			partial_clause[9][161] 	= partial_clause_prev[9][161] & 1'b1;
			partial_clause[9][162] 	= partial_clause_prev[9][162] & 1'b1;
			partial_clause[9][163] 	= partial_clause_prev[9][163] & 1'b1;
			partial_clause[9][164] 	= partial_clause_prev[9][164] & 1'b1;
			partial_clause[9][165] 	= partial_clause_prev[9][165] & ~x[52] & ~x[53];
			partial_clause[9][166] 	= partial_clause_prev[9][166] & 1'b1;
			partial_clause[9][167] 	= partial_clause_prev[9][167] & ~x[19] & ~x[47];
			partial_clause[9][168] 	= partial_clause_prev[9][168] & 1'b1;
			partial_clause[9][169] 	= partial_clause_prev[9][169] & 1'b1;
			partial_clause[9][170] 	= partial_clause_prev[9][170] & ~x[52];
			partial_clause[9][171] 	= partial_clause_prev[9][171] & 1'b1;
			partial_clause[9][172] 	= partial_clause_prev[9][172] & ~x[17];
			partial_clause[9][173] 	= partial_clause_prev[9][173] & 1'b1;
			partial_clause[9][174] 	= partial_clause_prev[9][174] & 1'b1;
			partial_clause[9][175] 	= partial_clause_prev[9][175] & 1'b1;
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & 1'b1;
			partial_clause[9][178] 	= partial_clause_prev[9][178] & 1'b1;
			partial_clause[9][179] 	= partial_clause_prev[9][179] & 1'b1;
			partial_clause[9][180] 	= partial_clause_prev[9][180] & 1'b1;
			partial_clause[9][181] 	= partial_clause_prev[9][181] & 1'b1;
			partial_clause[9][182] 	= partial_clause_prev[9][182] & ~x[18] & ~x[45];
			partial_clause[9][183] 	= partial_clause_prev[9][183] & 1'b1;
			partial_clause[9][184] 	= partial_clause_prev[9][184] & 1'b1;
			partial_clause[9][185] 	= partial_clause_prev[9][185] & 1'b1;
			partial_clause[9][186] 	= partial_clause_prev[9][186] & 1'b1;
			partial_clause[9][187] 	= partial_clause_prev[9][187] & 1'b1;
			partial_clause[9][188] 	= partial_clause_prev[9][188] & 1'b1;
			partial_clause[9][189] 	= partial_clause_prev[9][189] & ~x[15];
			partial_clause[9][190] 	= partial_clause_prev[9][190] & 1'b1;
			partial_clause[9][191] 	= partial_clause_prev[9][191] & 1'b1;
			partial_clause[9][192] 	= partial_clause_prev[9][192] & 1'b1;
			partial_clause[9][193] 	= partial_clause_prev[9][193] & 1'b1;
			partial_clause[9][194] 	= partial_clause_prev[9][194] & 1'b1;
			partial_clause[9][195] 	= partial_clause_prev[9][195] & 1'b1;
			partial_clause[9][196] 	= partial_clause_prev[9][196] & ~x[17];
			partial_clause[9][197] 	= partial_clause_prev[9][197] & 1'b1;
			partial_clause[9][198] 	= partial_clause_prev[9][198] & 1'b1;
			partial_clause[9][199] 	= partial_clause_prev[9][199] & x[59];
		end
	end
endmodule


module HCB_7 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & ~x[14];
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & ~x[43];
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & x[26];
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & ~x[15];
			partial_clause[0][11] 	= partial_clause_prev[0][11] & ~x[42];
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & ~x[15] & ~x[43];
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & x[45] & ~x[49];
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & x[8];
			partial_clause[0][18] 	= partial_clause_prev[0][18] & ~x[41];
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & x[38];
			partial_clause[0][24] 	= partial_clause_prev[0][24] & x[8] & ~x[22];
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & x[10];
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & ~x[40];
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & x[34];
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & x[9];
			partial_clause[0][45] 	= partial_clause_prev[0][45] & x[27];
			partial_clause[0][46] 	= partial_clause_prev[0][46] & ~x[16] & ~x[44];
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & ~x[13];
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & x[56];
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & x[20];
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & x[24];
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & ~x[14];
			partial_clause[0][64] 	= partial_clause_prev[0][64] & ~x[16] & ~x[43];
			partial_clause[0][65] 	= partial_clause_prev[0][65] & ~x[42];
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & ~x[16];
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & ~x[14] & x[38];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & ~x[42];
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & ~x[43];
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & ~x[40];
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & x[37];
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & x[33];
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & x[17];
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & ~x[62];
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			partial_clause[0][100] 	= partial_clause_prev[0][100] & 1'b1;
			partial_clause[0][101] 	= partial_clause_prev[0][101] & x[14];
			partial_clause[0][102] 	= partial_clause_prev[0][102] & x[16];
			partial_clause[0][103] 	= partial_clause_prev[0][103] & 1'b1;
			partial_clause[0][104] 	= partial_clause_prev[0][104] & ~x[29];
			partial_clause[0][105] 	= partial_clause_prev[0][105] & 1'b1;
			partial_clause[0][106] 	= partial_clause_prev[0][106] & 1'b1;
			partial_clause[0][107] 	= partial_clause_prev[0][107] & 1'b1;
			partial_clause[0][108] 	= partial_clause_prev[0][108] & 1'b1;
			partial_clause[0][109] 	= partial_clause_prev[0][109] & 1'b1;
			partial_clause[0][110] 	= partial_clause_prev[0][110] & 1'b1;
			partial_clause[0][111] 	= partial_clause_prev[0][111] & x[15];
			partial_clause[0][112] 	= partial_clause_prev[0][112] & 1'b1;
			partial_clause[0][113] 	= partial_clause_prev[0][113] & 1'b1;
			partial_clause[0][114] 	= partial_clause_prev[0][114] & 1'b1;
			partial_clause[0][115] 	= partial_clause_prev[0][115] & 1'b1;
			partial_clause[0][116] 	= partial_clause_prev[0][116] & x[42];
			partial_clause[0][117] 	= partial_clause_prev[0][117] & 1'b1;
			partial_clause[0][118] 	= partial_clause_prev[0][118] & 1'b1;
			partial_clause[0][119] 	= partial_clause_prev[0][119] & 1'b1;
			partial_clause[0][120] 	= partial_clause_prev[0][120] & 1'b1;
			partial_clause[0][121] 	= partial_clause_prev[0][121] & 1'b1;
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & ~x[5] & ~x[7] & ~x[8];
			partial_clause[0][124] 	= partial_clause_prev[0][124] & 1'b1;
			partial_clause[0][125] 	= partial_clause_prev[0][125] & 1'b1;
			partial_clause[0][126] 	= partial_clause_prev[0][126] & 1'b1;
			partial_clause[0][127] 	= partial_clause_prev[0][127] & 1'b1;
			partial_clause[0][128] 	= partial_clause_prev[0][128] & ~x[51] & ~x[62];
			partial_clause[0][129] 	= partial_clause_prev[0][129] & 1'b1;
			partial_clause[0][130] 	= partial_clause_prev[0][130] & ~x[36] & ~x[61] & ~x[63];
			partial_clause[0][131] 	= partial_clause_prev[0][131] & 1'b1;
			partial_clause[0][132] 	= partial_clause_prev[0][132] & 1'b1;
			partial_clause[0][133] 	= partial_clause_prev[0][133] & 1'b1;
			partial_clause[0][134] 	= partial_clause_prev[0][134] & 1'b1;
			partial_clause[0][135] 	= partial_clause_prev[0][135] & 1'b1;
			partial_clause[0][136] 	= partial_clause_prev[0][136] & ~x[9] & ~x[10];
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & 1'b1;
			partial_clause[0][139] 	= partial_clause_prev[0][139] & 1'b1;
			partial_clause[0][140] 	= partial_clause_prev[0][140] & 1'b1;
			partial_clause[0][141] 	= partial_clause_prev[0][141] & 1'b1;
			partial_clause[0][142] 	= partial_clause_prev[0][142] & ~x[35];
			partial_clause[0][143] 	= partial_clause_prev[0][143] & 1'b1;
			partial_clause[0][144] 	= partial_clause_prev[0][144] & 1'b1;
			partial_clause[0][145] 	= partial_clause_prev[0][145] & ~x[5] & ~x[36] & ~x[38];
			partial_clause[0][146] 	= partial_clause_prev[0][146] & 1'b1;
			partial_clause[0][147] 	= partial_clause_prev[0][147] & 1'b1;
			partial_clause[0][148] 	= partial_clause_prev[0][148] & 1'b1;
			partial_clause[0][149] 	= partial_clause_prev[0][149] & 1'b1;
			partial_clause[0][150] 	= partial_clause_prev[0][150] & x[14];
			partial_clause[0][151] 	= partial_clause_prev[0][151] & 1'b1;
			partial_clause[0][152] 	= partial_clause_prev[0][152] & 1'b1;
			partial_clause[0][153] 	= partial_clause_prev[0][153] & 1'b1;
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & 1'b1;
			partial_clause[0][156] 	= partial_clause_prev[0][156] & 1'b1;
			partial_clause[0][157] 	= partial_clause_prev[0][157] & x[12];
			partial_clause[0][158] 	= partial_clause_prev[0][158] & 1'b1;
			partial_clause[0][159] 	= partial_clause_prev[0][159] & x[41];
			partial_clause[0][160] 	= partial_clause_prev[0][160] & 1'b1;
			partial_clause[0][161] 	= partial_clause_prev[0][161] & 1'b1;
			partial_clause[0][162] 	= partial_clause_prev[0][162] & 1'b1;
			partial_clause[0][163] 	= partial_clause_prev[0][163] & 1'b1;
			partial_clause[0][164] 	= partial_clause_prev[0][164] & ~x[8] & ~x[38];
			partial_clause[0][165] 	= partial_clause_prev[0][165] & ~x[24];
			partial_clause[0][166] 	= partial_clause_prev[0][166] & x[14];
			partial_clause[0][167] 	= partial_clause_prev[0][167] & 1'b1;
			partial_clause[0][168] 	= partial_clause_prev[0][168] & 1'b1;
			partial_clause[0][169] 	= partial_clause_prev[0][169] & 1'b1;
			partial_clause[0][170] 	= partial_clause_prev[0][170] & 1'b1;
			partial_clause[0][171] 	= partial_clause_prev[0][171] & 1'b1;
			partial_clause[0][172] 	= partial_clause_prev[0][172] & 1'b1;
			partial_clause[0][173] 	= partial_clause_prev[0][173] & 1'b1;
			partial_clause[0][174] 	= partial_clause_prev[0][174] & 1'b1;
			partial_clause[0][175] 	= partial_clause_prev[0][175] & 1'b1;
			partial_clause[0][176] 	= partial_clause_prev[0][176] & 1'b1;
			partial_clause[0][177] 	= partial_clause_prev[0][177] & 1'b1;
			partial_clause[0][178] 	= partial_clause_prev[0][178] & 1'b1;
			partial_clause[0][179] 	= partial_clause_prev[0][179] & 1'b1;
			partial_clause[0][180] 	= partial_clause_prev[0][180] & 1'b1;
			partial_clause[0][181] 	= partial_clause_prev[0][181] & 1'b1;
			partial_clause[0][182] 	= partial_clause_prev[0][182] & 1'b1;
			partial_clause[0][183] 	= partial_clause_prev[0][183] & ~x[7] & ~x[38];
			partial_clause[0][184] 	= partial_clause_prev[0][184] & ~x[63];
			partial_clause[0][185] 	= partial_clause_prev[0][185] & 1'b1;
			partial_clause[0][186] 	= partial_clause_prev[0][186] & 1'b1;
			partial_clause[0][187] 	= partial_clause_prev[0][187] & 1'b1;
			partial_clause[0][188] 	= partial_clause_prev[0][188] & 1'b1;
			partial_clause[0][189] 	= partial_clause_prev[0][189] & x[42];
			partial_clause[0][190] 	= partial_clause_prev[0][190] & 1'b1;
			partial_clause[0][191] 	= partial_clause_prev[0][191] & 1'b1;
			partial_clause[0][192] 	= partial_clause_prev[0][192] & 1'b1;
			partial_clause[0][193] 	= partial_clause_prev[0][193] & 1'b1;
			partial_clause[0][194] 	= partial_clause_prev[0][194] & x[13] & x[14];
			partial_clause[0][195] 	= partial_clause_prev[0][195] & 1'b1;
			partial_clause[0][196] 	= partial_clause_prev[0][196] & 1'b1;
			partial_clause[0][197] 	= partial_clause_prev[0][197] & 1'b1;
			partial_clause[0][198] 	= partial_clause_prev[0][198] & 1'b1;
			partial_clause[0][199] 	= partial_clause_prev[0][199] & x[13] & x[14];
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[21] & x[40];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & ~x[16];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & ~x[39];
			partial_clause[1][9] 	= partial_clause_prev[1][9] & ~x[45];
			partial_clause[1][10] 	= partial_clause_prev[1][10] & ~x[39] & x[42];
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & ~x[39];
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & ~x[46];
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & ~x[11] & x[14];
			partial_clause[1][30] 	= partial_clause_prev[1][30] & x[25];
			partial_clause[1][31] 	= partial_clause_prev[1][31] & x[57];
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & ~x[44];
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & x[13];
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & ~x[10];
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & x[13];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & x[42];
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & ~x[7];
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & ~x[17];
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & x[58];
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & x[13] & ~x[45];
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & x[41];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & ~x[39];
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & x[42];
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & ~x[39];
			partial_clause[1][90] 	= partial_clause_prev[1][90] & ~x[16];
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			partial_clause[1][100] 	= partial_clause_prev[1][100] & x[46];
			partial_clause[1][101] 	= partial_clause_prev[1][101] & 1'b1;
			partial_clause[1][102] 	= partial_clause_prev[1][102] & 1'b1;
			partial_clause[1][103] 	= partial_clause_prev[1][103] & x[62];
			partial_clause[1][104] 	= partial_clause_prev[1][104] & 1'b1;
			partial_clause[1][105] 	= partial_clause_prev[1][105] & 1'b1;
			partial_clause[1][106] 	= partial_clause_prev[1][106] & 1'b1;
			partial_clause[1][107] 	= partial_clause_prev[1][107] & 1'b1;
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & 1'b1;
			partial_clause[1][110] 	= partial_clause_prev[1][110] & 1'b1;
			partial_clause[1][111] 	= partial_clause_prev[1][111] & 1'b1;
			partial_clause[1][112] 	= partial_clause_prev[1][112] & 1'b1;
			partial_clause[1][113] 	= partial_clause_prev[1][113] & x[47];
			partial_clause[1][114] 	= partial_clause_prev[1][114] & x[10];
			partial_clause[1][115] 	= partial_clause_prev[1][115] & 1'b1;
			partial_clause[1][116] 	= partial_clause_prev[1][116] & 1'b1;
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & 1'b1;
			partial_clause[1][119] 	= partial_clause_prev[1][119] & 1'b1;
			partial_clause[1][120] 	= partial_clause_prev[1][120] & 1'b1;
			partial_clause[1][121] 	= partial_clause_prev[1][121] & x[49];
			partial_clause[1][122] 	= partial_clause_prev[1][122] & 1'b1;
			partial_clause[1][123] 	= partial_clause_prev[1][123] & 1'b1;
			partial_clause[1][124] 	= partial_clause_prev[1][124] & 1'b1;
			partial_clause[1][125] 	= partial_clause_prev[1][125] & 1'b1;
			partial_clause[1][126] 	= partial_clause_prev[1][126] & 1'b1;
			partial_clause[1][127] 	= partial_clause_prev[1][127] & ~x[57];
			partial_clause[1][128] 	= partial_clause_prev[1][128] & 1'b1;
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & 1'b1;
			partial_clause[1][131] 	= partial_clause_prev[1][131] & x[63];
			partial_clause[1][132] 	= partial_clause_prev[1][132] & 1'b1;
			partial_clause[1][133] 	= partial_clause_prev[1][133] & x[63];
			partial_clause[1][134] 	= partial_clause_prev[1][134] & 1'b1;
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & 1'b1;
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & 1'b1;
			partial_clause[1][139] 	= partial_clause_prev[1][139] & 1'b1;
			partial_clause[1][140] 	= partial_clause_prev[1][140] & 1'b1;
			partial_clause[1][141] 	= partial_clause_prev[1][141] & 1'b1;
			partial_clause[1][142] 	= partial_clause_prev[1][142] & 1'b1;
			partial_clause[1][143] 	= partial_clause_prev[1][143] & 1'b1;
			partial_clause[1][144] 	= partial_clause_prev[1][144] & 1'b1;
			partial_clause[1][145] 	= partial_clause_prev[1][145] & 1'b1;
			partial_clause[1][146] 	= partial_clause_prev[1][146] & 1'b1;
			partial_clause[1][147] 	= partial_clause_prev[1][147] & 1'b1;
			partial_clause[1][148] 	= partial_clause_prev[1][148] & 1'b1;
			partial_clause[1][149] 	= partial_clause_prev[1][149] & x[37];
			partial_clause[1][150] 	= partial_clause_prev[1][150] & ~x[13] & ~x[14];
			partial_clause[1][151] 	= partial_clause_prev[1][151] & 1'b1;
			partial_clause[1][152] 	= partial_clause_prev[1][152] & 1'b1;
			partial_clause[1][153] 	= partial_clause_prev[1][153] & 1'b1;
			partial_clause[1][154] 	= partial_clause_prev[1][154] & 1'b1;
			partial_clause[1][155] 	= partial_clause_prev[1][155] & 1'b1;
			partial_clause[1][156] 	= partial_clause_prev[1][156] & 1'b1;
			partial_clause[1][157] 	= partial_clause_prev[1][157] & ~x[42];
			partial_clause[1][158] 	= partial_clause_prev[1][158] & 1'b1;
			partial_clause[1][159] 	= partial_clause_prev[1][159] & 1'b1;
			partial_clause[1][160] 	= partial_clause_prev[1][160] & 1'b1;
			partial_clause[1][161] 	= partial_clause_prev[1][161] & x[8];
			partial_clause[1][162] 	= partial_clause_prev[1][162] & 1'b1;
			partial_clause[1][163] 	= partial_clause_prev[1][163] & 1'b1;
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & 1'b1;
			partial_clause[1][166] 	= partial_clause_prev[1][166] & 1'b1;
			partial_clause[1][167] 	= partial_clause_prev[1][167] & 1'b1;
			partial_clause[1][168] 	= partial_clause_prev[1][168] & 1'b1;
			partial_clause[1][169] 	= partial_clause_prev[1][169] & 1'b1;
			partial_clause[1][170] 	= partial_clause_prev[1][170] & 1'b1;
			partial_clause[1][171] 	= partial_clause_prev[1][171] & 1'b1;
			partial_clause[1][172] 	= partial_clause_prev[1][172] & 1'b1;
			partial_clause[1][173] 	= partial_clause_prev[1][173] & 1'b1;
			partial_clause[1][174] 	= partial_clause_prev[1][174] & 1'b1;
			partial_clause[1][175] 	= partial_clause_prev[1][175] & 1'b1;
			partial_clause[1][176] 	= partial_clause_prev[1][176] & x[17] & ~x[43];
			partial_clause[1][177] 	= partial_clause_prev[1][177] & 1'b1;
			partial_clause[1][178] 	= partial_clause_prev[1][178] & 1'b1;
			partial_clause[1][179] 	= partial_clause_prev[1][179] & 1'b1;
			partial_clause[1][180] 	= partial_clause_prev[1][180] & 1'b1;
			partial_clause[1][181] 	= partial_clause_prev[1][181] & 1'b1;
			partial_clause[1][182] 	= partial_clause_prev[1][182] & 1'b1;
			partial_clause[1][183] 	= partial_clause_prev[1][183] & x[35];
			partial_clause[1][184] 	= partial_clause_prev[1][184] & 1'b1;
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & 1'b1;
			partial_clause[1][187] 	= partial_clause_prev[1][187] & 1'b1;
			partial_clause[1][188] 	= partial_clause_prev[1][188] & 1'b1;
			partial_clause[1][189] 	= partial_clause_prev[1][189] & ~x[15];
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & x[18];
			partial_clause[1][192] 	= partial_clause_prev[1][192] & 1'b1;
			partial_clause[1][193] 	= partial_clause_prev[1][193] & ~x[31];
			partial_clause[1][194] 	= partial_clause_prev[1][194] & ~x[41];
			partial_clause[1][195] 	= partial_clause_prev[1][195] & 1'b1;
			partial_clause[1][196] 	= partial_clause_prev[1][196] & 1'b1;
			partial_clause[1][197] 	= partial_clause_prev[1][197] & 1'b1;
			partial_clause[1][198] 	= partial_clause_prev[1][198] & x[17];
			partial_clause[1][199] 	= partial_clause_prev[1][199] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & x[53];
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & x[25];
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & x[33];
			partial_clause[2][22] 	= partial_clause_prev[2][22] & x[44] & x[46];
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & x[15];
			partial_clause[2][27] 	= partial_clause_prev[2][27] & ~x[48];
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & x[59];
			partial_clause[2][37] 	= partial_clause_prev[2][37] & x[43];
			partial_clause[2][38] 	= partial_clause_prev[2][38] & ~x[5];
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & ~x[48] & ~x[49];
			partial_clause[2][43] 	= partial_clause_prev[2][43] & x[52];
			partial_clause[2][44] 	= partial_clause_prev[2][44] & x[41] & ~x[46];
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & x[53];
			partial_clause[2][47] 	= partial_clause_prev[2][47] & ~x[47] & ~x[48];
			partial_clause[2][48] 	= partial_clause_prev[2][48] & x[53];
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & x[35];
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & x[25];
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & x[17];
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & x[45];
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & x[43];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & x[25];
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & x[26];
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & x[11];
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & x[7];
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & x[61];
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & x[53];
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & x[53];
			partial_clause[2][93] 	= partial_clause_prev[2][93] & ~x[20];
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & ~x[48] & ~x[50];
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & x[45] & x[49];
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			partial_clause[2][100] 	= partial_clause_prev[2][100] & ~x[25] & ~x[52];
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & ~x[10];
			partial_clause[2][103] 	= partial_clause_prev[2][103] & 1'b1;
			partial_clause[2][104] 	= partial_clause_prev[2][104] & ~x[19] & ~x[46];
			partial_clause[2][105] 	= partial_clause_prev[2][105] & 1'b1;
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & 1'b1;
			partial_clause[2][108] 	= partial_clause_prev[2][108] & 1'b1;
			partial_clause[2][109] 	= partial_clause_prev[2][109] & 1'b1;
			partial_clause[2][110] 	= partial_clause_prev[2][110] & 1'b1;
			partial_clause[2][111] 	= partial_clause_prev[2][111] & 1'b1;
			partial_clause[2][112] 	= partial_clause_prev[2][112] & 1'b1;
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & ~x[5];
			partial_clause[2][115] 	= partial_clause_prev[2][115] & 1'b1;
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & 1'b1;
			partial_clause[2][118] 	= partial_clause_prev[2][118] & 1'b1;
			partial_clause[2][119] 	= partial_clause_prev[2][119] & 1'b1;
			partial_clause[2][120] 	= partial_clause_prev[2][120] & 1'b1;
			partial_clause[2][121] 	= partial_clause_prev[2][121] & ~x[63];
			partial_clause[2][122] 	= partial_clause_prev[2][122] & 1'b1;
			partial_clause[2][123] 	= partial_clause_prev[2][123] & 1'b1;
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & ~x[11] & ~x[12] & ~x[40] & ~x[44];
			partial_clause[2][126] 	= partial_clause_prev[2][126] & 1'b1;
			partial_clause[2][127] 	= partial_clause_prev[2][127] & 1'b1;
			partial_clause[2][128] 	= partial_clause_prev[2][128] & 1'b1;
			partial_clause[2][129] 	= partial_clause_prev[2][129] & 1'b1;
			partial_clause[2][130] 	= partial_clause_prev[2][130] & 1'b1;
			partial_clause[2][131] 	= partial_clause_prev[2][131] & ~x[10];
			partial_clause[2][132] 	= partial_clause_prev[2][132] & 1'b1;
			partial_clause[2][133] 	= partial_clause_prev[2][133] & 1'b1;
			partial_clause[2][134] 	= partial_clause_prev[2][134] & 1'b1;
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & 1'b1;
			partial_clause[2][137] 	= partial_clause_prev[2][137] & x[8];
			partial_clause[2][138] 	= partial_clause_prev[2][138] & 1'b1;
			partial_clause[2][139] 	= partial_clause_prev[2][139] & 1'b1;
			partial_clause[2][140] 	= partial_clause_prev[2][140] & 1'b1;
			partial_clause[2][141] 	= partial_clause_prev[2][141] & 1'b1;
			partial_clause[2][142] 	= partial_clause_prev[2][142] & 1'b1;
			partial_clause[2][143] 	= partial_clause_prev[2][143] & 1'b1;
			partial_clause[2][144] 	= partial_clause_prev[2][144] & 1'b1;
			partial_clause[2][145] 	= partial_clause_prev[2][145] & 1'b1;
			partial_clause[2][146] 	= partial_clause_prev[2][146] & ~x[5] & ~x[6] & ~x[7];
			partial_clause[2][147] 	= partial_clause_prev[2][147] & 1'b1;
			partial_clause[2][148] 	= partial_clause_prev[2][148] & ~x[8] & ~x[25] & ~x[38];
			partial_clause[2][149] 	= partial_clause_prev[2][149] & ~x[23];
			partial_clause[2][150] 	= partial_clause_prev[2][150] & ~x[39];
			partial_clause[2][151] 	= partial_clause_prev[2][151] & 1'b1;
			partial_clause[2][152] 	= partial_clause_prev[2][152] & 1'b1;
			partial_clause[2][153] 	= partial_clause_prev[2][153] & 1'b1;
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & ~x[21];
			partial_clause[2][156] 	= partial_clause_prev[2][156] & 1'b1;
			partial_clause[2][157] 	= partial_clause_prev[2][157] & 1'b1;
			partial_clause[2][158] 	= partial_clause_prev[2][158] & 1'b1;
			partial_clause[2][159] 	= partial_clause_prev[2][159] & 1'b1;
			partial_clause[2][160] 	= partial_clause_prev[2][160] & 1'b1;
			partial_clause[2][161] 	= partial_clause_prev[2][161] & ~x[19] & ~x[36];
			partial_clause[2][162] 	= partial_clause_prev[2][162] & ~x[7];
			partial_clause[2][163] 	= partial_clause_prev[2][163] & 1'b1;
			partial_clause[2][164] 	= partial_clause_prev[2][164] & 1'b1;
			partial_clause[2][165] 	= partial_clause_prev[2][165] & 1'b1;
			partial_clause[2][166] 	= partial_clause_prev[2][166] & ~x[40];
			partial_clause[2][167] 	= partial_clause_prev[2][167] & x[8];
			partial_clause[2][168] 	= partial_clause_prev[2][168] & ~x[34];
			partial_clause[2][169] 	= partial_clause_prev[2][169] & ~x[21] & ~x[49];
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & 1'b1;
			partial_clause[2][173] 	= partial_clause_prev[2][173] & 1'b1;
			partial_clause[2][174] 	= partial_clause_prev[2][174] & 1'b1;
			partial_clause[2][175] 	= partial_clause_prev[2][175] & 1'b1;
			partial_clause[2][176] 	= partial_clause_prev[2][176] & 1'b1;
			partial_clause[2][177] 	= partial_clause_prev[2][177] & 1'b1;
			partial_clause[2][178] 	= partial_clause_prev[2][178] & 1'b1;
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & 1'b1;
			partial_clause[2][181] 	= partial_clause_prev[2][181] & ~x[22];
			partial_clause[2][182] 	= partial_clause_prev[2][182] & 1'b1;
			partial_clause[2][183] 	= partial_clause_prev[2][183] & 1'b1;
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & 1'b1;
			partial_clause[2][186] 	= partial_clause_prev[2][186] & 1'b1;
			partial_clause[2][187] 	= partial_clause_prev[2][187] & 1'b1;
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & ~x[8];
			partial_clause[2][190] 	= partial_clause_prev[2][190] & ~x[39];
			partial_clause[2][191] 	= partial_clause_prev[2][191] & 1'b1;
			partial_clause[2][192] 	= partial_clause_prev[2][192] & 1'b1;
			partial_clause[2][193] 	= partial_clause_prev[2][193] & 1'b1;
			partial_clause[2][194] 	= partial_clause_prev[2][194] & 1'b1;
			partial_clause[2][195] 	= partial_clause_prev[2][195] & 1'b1;
			partial_clause[2][196] 	= partial_clause_prev[2][196] & 1'b1;
			partial_clause[2][197] 	= partial_clause_prev[2][197] & 1'b1;
			partial_clause[2][198] 	= partial_clause_prev[2][198] & ~x[23] & ~x[36];
			partial_clause[2][199] 	= partial_clause_prev[2][199] & ~x[7] & ~x[36] & ~x[38];
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & ~x[37] & ~x[38] & ~x[39] & ~x[40];
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & ~x[11] & ~x[42];
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & x[26];
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & ~x[10];
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & ~x[36];
			partial_clause[3][25] 	= partial_clause_prev[3][25] & x[60];
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & ~x[38] & ~x[39];
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & ~x[37];
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & ~x[37] & ~x[38];
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & ~x[8] & ~x[39] & ~x[40];
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & ~x[39];
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & x[48];
			partial_clause[3][58] 	= partial_clause_prev[3][58] & ~x[8] & ~x[38];
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & ~x[38];
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & 1'b1;
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & x[54];
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & x[60];
			partial_clause[3][71] 	= partial_clause_prev[3][71] & ~x[41];
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & x[29];
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & ~x[12] & ~x[14];
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & x[31];
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & x[18];
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & ~x[14];
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			partial_clause[3][100] 	= partial_clause_prev[3][100] & x[44];
			partial_clause[3][101] 	= partial_clause_prev[3][101] & 1'b1;
			partial_clause[3][102] 	= partial_clause_prev[3][102] & x[14] & ~x[18] & ~x[45];
			partial_clause[3][103] 	= partial_clause_prev[3][103] & 1'b1;
			partial_clause[3][104] 	= partial_clause_prev[3][104] & 1'b1;
			partial_clause[3][105] 	= partial_clause_prev[3][105] & 1'b1;
			partial_clause[3][106] 	= partial_clause_prev[3][106] & ~x[45];
			partial_clause[3][107] 	= partial_clause_prev[3][107] & 1'b1;
			partial_clause[3][108] 	= partial_clause_prev[3][108] & x[11] & x[38];
			partial_clause[3][109] 	= partial_clause_prev[3][109] & 1'b1;
			partial_clause[3][110] 	= partial_clause_prev[3][110] & x[43];
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & 1'b1;
			partial_clause[3][113] 	= partial_clause_prev[3][113] & 1'b1;
			partial_clause[3][114] 	= partial_clause_prev[3][114] & x[37];
			partial_clause[3][115] 	= partial_clause_prev[3][115] & 1'b1;
			partial_clause[3][116] 	= partial_clause_prev[3][116] & 1'b1;
			partial_clause[3][117] 	= partial_clause_prev[3][117] & 1'b1;
			partial_clause[3][118] 	= partial_clause_prev[3][118] & ~x[21] & ~x[46] & ~x[47];
			partial_clause[3][119] 	= partial_clause_prev[3][119] & 1'b1;
			partial_clause[3][120] 	= partial_clause_prev[3][120] & 1'b1;
			partial_clause[3][121] 	= partial_clause_prev[3][121] & 1'b1;
			partial_clause[3][122] 	= partial_clause_prev[3][122] & 1'b1;
			partial_clause[3][123] 	= partial_clause_prev[3][123] & x[12];
			partial_clause[3][124] 	= partial_clause_prev[3][124] & x[12];
			partial_clause[3][125] 	= partial_clause_prev[3][125] & 1'b1;
			partial_clause[3][126] 	= partial_clause_prev[3][126] & 1'b1;
			partial_clause[3][127] 	= partial_clause_prev[3][127] & 1'b1;
			partial_clause[3][128] 	= partial_clause_prev[3][128] & 1'b1;
			partial_clause[3][129] 	= partial_clause_prev[3][129] & 1'b1;
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & 1'b1;
			partial_clause[3][132] 	= partial_clause_prev[3][132] & 1'b1;
			partial_clause[3][133] 	= partial_clause_prev[3][133] & 1'b1;
			partial_clause[3][134] 	= partial_clause_prev[3][134] & 1'b1;
			partial_clause[3][135] 	= partial_clause_prev[3][135] & 1'b1;
			partial_clause[3][136] 	= partial_clause_prev[3][136] & 1'b1;
			partial_clause[3][137] 	= partial_clause_prev[3][137] & 1'b1;
			partial_clause[3][138] 	= partial_clause_prev[3][138] & 1'b1;
			partial_clause[3][139] 	= partial_clause_prev[3][139] & x[44];
			partial_clause[3][140] 	= partial_clause_prev[3][140] & 1'b1;
			partial_clause[3][141] 	= partial_clause_prev[3][141] & 1'b1;
			partial_clause[3][142] 	= partial_clause_prev[3][142] & x[12] & x[39];
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & 1'b1;
			partial_clause[3][145] 	= partial_clause_prev[3][145] & ~x[45];
			partial_clause[3][146] 	= partial_clause_prev[3][146] & 1'b1;
			partial_clause[3][147] 	= partial_clause_prev[3][147] & 1'b1;
			partial_clause[3][148] 	= partial_clause_prev[3][148] & 1'b1;
			partial_clause[3][149] 	= partial_clause_prev[3][149] & 1'b1;
			partial_clause[3][150] 	= partial_clause_prev[3][150] & 1'b1;
			partial_clause[3][151] 	= partial_clause_prev[3][151] & 1'b1;
			partial_clause[3][152] 	= partial_clause_prev[3][152] & 1'b1;
			partial_clause[3][153] 	= partial_clause_prev[3][153] & 1'b1;
			partial_clause[3][154] 	= partial_clause_prev[3][154] & 1'b1;
			partial_clause[3][155] 	= partial_clause_prev[3][155] & 1'b1;
			partial_clause[3][156] 	= partial_clause_prev[3][156] & x[14];
			partial_clause[3][157] 	= partial_clause_prev[3][157] & 1'b1;
			partial_clause[3][158] 	= partial_clause_prev[3][158] & 1'b1;
			partial_clause[3][159] 	= partial_clause_prev[3][159] & 1'b1;
			partial_clause[3][160] 	= partial_clause_prev[3][160] & 1'b1;
			partial_clause[3][161] 	= partial_clause_prev[3][161] & 1'b1;
			partial_clause[3][162] 	= partial_clause_prev[3][162] & 1'b1;
			partial_clause[3][163] 	= partial_clause_prev[3][163] & 1'b1;
			partial_clause[3][164] 	= partial_clause_prev[3][164] & 1'b1;
			partial_clause[3][165] 	= partial_clause_prev[3][165] & 1'b1;
			partial_clause[3][166] 	= partial_clause_prev[3][166] & x[38];
			partial_clause[3][167] 	= partial_clause_prev[3][167] & x[41];
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & 1'b1;
			partial_clause[3][170] 	= partial_clause_prev[3][170] & 1'b1;
			partial_clause[3][171] 	= partial_clause_prev[3][171] & ~x[20] & x[42];
			partial_clause[3][172] 	= partial_clause_prev[3][172] & 1'b1;
			partial_clause[3][173] 	= partial_clause_prev[3][173] & ~x[49];
			partial_clause[3][174] 	= partial_clause_prev[3][174] & x[37];
			partial_clause[3][175] 	= partial_clause_prev[3][175] & x[41];
			partial_clause[3][176] 	= partial_clause_prev[3][176] & 1'b1;
			partial_clause[3][177] 	= partial_clause_prev[3][177] & 1'b1;
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & 1'b1;
			partial_clause[3][180] 	= partial_clause_prev[3][180] & 1'b1;
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & 1'b1;
			partial_clause[3][183] 	= partial_clause_prev[3][183] & 1'b1;
			partial_clause[3][184] 	= partial_clause_prev[3][184] & 1'b1;
			partial_clause[3][185] 	= partial_clause_prev[3][185] & 1'b1;
			partial_clause[3][186] 	= partial_clause_prev[3][186] & 1'b1;
			partial_clause[3][187] 	= partial_clause_prev[3][187] & 1'b1;
			partial_clause[3][188] 	= partial_clause_prev[3][188] & 1'b1;
			partial_clause[3][189] 	= partial_clause_prev[3][189] & 1'b1;
			partial_clause[3][190] 	= partial_clause_prev[3][190] & 1'b1;
			partial_clause[3][191] 	= partial_clause_prev[3][191] & ~x[18];
			partial_clause[3][192] 	= partial_clause_prev[3][192] & 1'b1;
			partial_clause[3][193] 	= partial_clause_prev[3][193] & 1'b1;
			partial_clause[3][194] 	= partial_clause_prev[3][194] & 1'b1;
			partial_clause[3][195] 	= partial_clause_prev[3][195] & 1'b1;
			partial_clause[3][196] 	= partial_clause_prev[3][196] & 1'b1;
			partial_clause[3][197] 	= partial_clause_prev[3][197] & 1'b1;
			partial_clause[3][198] 	= partial_clause_prev[3][198] & ~x[18];
			partial_clause[3][199] 	= partial_clause_prev[3][199] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & x[13] & x[18];
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & 1'b1;
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & x[42];
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & x[27];
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & ~x[23];
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & 1'b1;
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & ~x[21];
			partial_clause[4][54] 	= partial_clause_prev[4][54] & x[15];
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & x[43];
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & x[7] & x[43];
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & x[16];
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & x[14];
			partial_clause[4][82] 	= partial_clause_prev[4][82] & ~x[23];
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & x[13] & x[14] & x[15];
			partial_clause[4][100] 	= partial_clause_prev[4][100] & 1'b1;
			partial_clause[4][101] 	= partial_clause_prev[4][101] & 1'b1;
			partial_clause[4][102] 	= partial_clause_prev[4][102] & 1'b1;
			partial_clause[4][103] 	= partial_clause_prev[4][103] & 1'b1;
			partial_clause[4][104] 	= partial_clause_prev[4][104] & 1'b1;
			partial_clause[4][105] 	= partial_clause_prev[4][105] & 1'b1;
			partial_clause[4][106] 	= partial_clause_prev[4][106] & 1'b1;
			partial_clause[4][107] 	= partial_clause_prev[4][107] & 1'b1;
			partial_clause[4][108] 	= partial_clause_prev[4][108] & ~x[8];
			partial_clause[4][109] 	= partial_clause_prev[4][109] & ~x[21];
			partial_clause[4][110] 	= partial_clause_prev[4][110] & 1'b1;
			partial_clause[4][111] 	= partial_clause_prev[4][111] & 1'b1;
			partial_clause[4][112] 	= partial_clause_prev[4][112] & 1'b1;
			partial_clause[4][113] 	= partial_clause_prev[4][113] & 1'b1;
			partial_clause[4][114] 	= partial_clause_prev[4][114] & 1'b1;
			partial_clause[4][115] 	= partial_clause_prev[4][115] & 1'b1;
			partial_clause[4][116] 	= partial_clause_prev[4][116] & 1'b1;
			partial_clause[4][117] 	= partial_clause_prev[4][117] & ~x[46];
			partial_clause[4][118] 	= partial_clause_prev[4][118] & 1'b1;
			partial_clause[4][119] 	= partial_clause_prev[4][119] & 1'b1;
			partial_clause[4][120] 	= partial_clause_prev[4][120] & 1'b1;
			partial_clause[4][121] 	= partial_clause_prev[4][121] & ~x[19];
			partial_clause[4][122] 	= partial_clause_prev[4][122] & 1'b1;
			partial_clause[4][123] 	= partial_clause_prev[4][123] & 1'b1;
			partial_clause[4][124] 	= partial_clause_prev[4][124] & 1'b1;
			partial_clause[4][125] 	= partial_clause_prev[4][125] & 1'b1;
			partial_clause[4][126] 	= partial_clause_prev[4][126] & 1'b1;
			partial_clause[4][127] 	= partial_clause_prev[4][127] & ~x[41];
			partial_clause[4][128] 	= partial_clause_prev[4][128] & 1'b1;
			partial_clause[4][129] 	= partial_clause_prev[4][129] & 1'b1;
			partial_clause[4][130] 	= partial_clause_prev[4][130] & ~x[7] & ~x[15];
			partial_clause[4][131] 	= partial_clause_prev[4][131] & 1'b1;
			partial_clause[4][132] 	= partial_clause_prev[4][132] & ~x[16];
			partial_clause[4][133] 	= partial_clause_prev[4][133] & 1'b1;
			partial_clause[4][134] 	= partial_clause_prev[4][134] & 1'b1;
			partial_clause[4][135] 	= partial_clause_prev[4][135] & ~x[8] & ~x[35];
			partial_clause[4][136] 	= partial_clause_prev[4][136] & 1'b1;
			partial_clause[4][137] 	= partial_clause_prev[4][137] & 1'b1;
			partial_clause[4][138] 	= partial_clause_prev[4][138] & 1'b1;
			partial_clause[4][139] 	= partial_clause_prev[4][139] & 1'b1;
			partial_clause[4][140] 	= partial_clause_prev[4][140] & ~x[35];
			partial_clause[4][141] 	= partial_clause_prev[4][141] & 1'b1;
			partial_clause[4][142] 	= partial_clause_prev[4][142] & 1'b1;
			partial_clause[4][143] 	= partial_clause_prev[4][143] & 1'b1;
			partial_clause[4][144] 	= partial_clause_prev[4][144] & 1'b1;
			partial_clause[4][145] 	= partial_clause_prev[4][145] & 1'b1;
			partial_clause[4][146] 	= partial_clause_prev[4][146] & 1'b1;
			partial_clause[4][147] 	= partial_clause_prev[4][147] & 1'b1;
			partial_clause[4][148] 	= partial_clause_prev[4][148] & 1'b1;
			partial_clause[4][149] 	= partial_clause_prev[4][149] & 1'b1;
			partial_clause[4][150] 	= partial_clause_prev[4][150] & ~x[37];
			partial_clause[4][151] 	= partial_clause_prev[4][151] & 1'b1;
			partial_clause[4][152] 	= partial_clause_prev[4][152] & 1'b1;
			partial_clause[4][153] 	= partial_clause_prev[4][153] & ~x[43];
			partial_clause[4][154] 	= partial_clause_prev[4][154] & ~x[44];
			partial_clause[4][155] 	= partial_clause_prev[4][155] & 1'b1;
			partial_clause[4][156] 	= partial_clause_prev[4][156] & 1'b1;
			partial_clause[4][157] 	= partial_clause_prev[4][157] & ~x[21];
			partial_clause[4][158] 	= partial_clause_prev[4][158] & 1'b1;
			partial_clause[4][159] 	= partial_clause_prev[4][159] & 1'b1;
			partial_clause[4][160] 	= partial_clause_prev[4][160] & 1'b1;
			partial_clause[4][161] 	= partial_clause_prev[4][161] & ~x[8] & ~x[35];
			partial_clause[4][162] 	= partial_clause_prev[4][162] & 1'b1;
			partial_clause[4][163] 	= partial_clause_prev[4][163] & 1'b1;
			partial_clause[4][164] 	= partial_clause_prev[4][164] & 1'b1;
			partial_clause[4][165] 	= partial_clause_prev[4][165] & 1'b1;
			partial_clause[4][166] 	= partial_clause_prev[4][166] & 1'b1;
			partial_clause[4][167] 	= partial_clause_prev[4][167] & 1'b1;
			partial_clause[4][168] 	= partial_clause_prev[4][168] & 1'b1;
			partial_clause[4][169] 	= partial_clause_prev[4][169] & 1'b1;
			partial_clause[4][170] 	= partial_clause_prev[4][170] & ~x[8];
			partial_clause[4][171] 	= partial_clause_prev[4][171] & ~x[17];
			partial_clause[4][172] 	= partial_clause_prev[4][172] & ~x[42];
			partial_clause[4][173] 	= partial_clause_prev[4][173] & 1'b1;
			partial_clause[4][174] 	= partial_clause_prev[4][174] & 1'b1;
			partial_clause[4][175] 	= partial_clause_prev[4][175] & 1'b1;
			partial_clause[4][176] 	= partial_clause_prev[4][176] & 1'b1;
			partial_clause[4][177] 	= partial_clause_prev[4][177] & ~x[43];
			partial_clause[4][178] 	= partial_clause_prev[4][178] & 1'b1;
			partial_clause[4][179] 	= partial_clause_prev[4][179] & 1'b1;
			partial_clause[4][180] 	= partial_clause_prev[4][180] & 1'b1;
			partial_clause[4][181] 	= partial_clause_prev[4][181] & 1'b1;
			partial_clause[4][182] 	= partial_clause_prev[4][182] & 1'b1;
			partial_clause[4][183] 	= partial_clause_prev[4][183] & 1'b1;
			partial_clause[4][184] 	= partial_clause_prev[4][184] & 1'b1;
			partial_clause[4][185] 	= partial_clause_prev[4][185] & 1'b1;
			partial_clause[4][186] 	= partial_clause_prev[4][186] & 1'b1;
			partial_clause[4][187] 	= partial_clause_prev[4][187] & 1'b1;
			partial_clause[4][188] 	= partial_clause_prev[4][188] & 1'b1;
			partial_clause[4][189] 	= partial_clause_prev[4][189] & ~x[19];
			partial_clause[4][190] 	= partial_clause_prev[4][190] & 1'b1;
			partial_clause[4][191] 	= partial_clause_prev[4][191] & ~x[15];
			partial_clause[4][192] 	= partial_clause_prev[4][192] & 1'b1;
			partial_clause[4][193] 	= partial_clause_prev[4][193] & ~x[14];
			partial_clause[4][194] 	= partial_clause_prev[4][194] & 1'b1;
			partial_clause[4][195] 	= partial_clause_prev[4][195] & 1'b1;
			partial_clause[4][196] 	= partial_clause_prev[4][196] & 1'b1;
			partial_clause[4][197] 	= partial_clause_prev[4][197] & 1'b1;
			partial_clause[4][198] 	= partial_clause_prev[4][198] & 1'b1;
			partial_clause[4][199] 	= partial_clause_prev[4][199] & ~x[34];
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & ~x[7] & ~x[37];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & x[58];
			partial_clause[5][28] 	= partial_clause_prev[5][28] & ~x[38] & ~x[42];
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & ~x[36] & ~x[40];
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & ~x[35];
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & ~x[38] & ~x[43];
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & ~x[37] & ~x[40];
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & ~x[38];
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & x[51];
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & ~x[35];
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			partial_clause[5][100] 	= partial_clause_prev[5][100] & 1'b1;
			partial_clause[5][101] 	= partial_clause_prev[5][101] & 1'b1;
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & 1'b1;
			partial_clause[5][104] 	= partial_clause_prev[5][104] & 1'b1;
			partial_clause[5][105] 	= partial_clause_prev[5][105] & 1'b1;
			partial_clause[5][106] 	= partial_clause_prev[5][106] & 1'b1;
			partial_clause[5][107] 	= partial_clause_prev[5][107] & x[10];
			partial_clause[5][108] 	= partial_clause_prev[5][108] & 1'b1;
			partial_clause[5][109] 	= partial_clause_prev[5][109] & 1'b1;
			partial_clause[5][110] 	= partial_clause_prev[5][110] & 1'b1;
			partial_clause[5][111] 	= partial_clause_prev[5][111] & 1'b1;
			partial_clause[5][112] 	= partial_clause_prev[5][112] & 1'b1;
			partial_clause[5][113] 	= partial_clause_prev[5][113] & 1'b1;
			partial_clause[5][114] 	= partial_clause_prev[5][114] & 1'b1;
			partial_clause[5][115] 	= partial_clause_prev[5][115] & 1'b1;
			partial_clause[5][116] 	= partial_clause_prev[5][116] & 1'b1;
			partial_clause[5][117] 	= partial_clause_prev[5][117] & 1'b1;
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & 1'b1;
			partial_clause[5][120] 	= partial_clause_prev[5][120] & 1'b1;
			partial_clause[5][121] 	= partial_clause_prev[5][121] & 1'b1;
			partial_clause[5][122] 	= partial_clause_prev[5][122] & x[14];
			partial_clause[5][123] 	= partial_clause_prev[5][123] & 1'b1;
			partial_clause[5][124] 	= partial_clause_prev[5][124] & 1'b1;
			partial_clause[5][125] 	= partial_clause_prev[5][125] & ~x[34];
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & ~x[21] & ~x[35];
			partial_clause[5][128] 	= partial_clause_prev[5][128] & x[12];
			partial_clause[5][129] 	= partial_clause_prev[5][129] & 1'b1;
			partial_clause[5][130] 	= partial_clause_prev[5][130] & 1'b1;
			partial_clause[5][131] 	= partial_clause_prev[5][131] & x[42];
			partial_clause[5][132] 	= partial_clause_prev[5][132] & ~x[63];
			partial_clause[5][133] 	= partial_clause_prev[5][133] & 1'b1;
			partial_clause[5][134] 	= partial_clause_prev[5][134] & x[10];
			partial_clause[5][135] 	= partial_clause_prev[5][135] & 1'b1;
			partial_clause[5][136] 	= partial_clause_prev[5][136] & 1'b1;
			partial_clause[5][137] 	= partial_clause_prev[5][137] & 1'b1;
			partial_clause[5][138] 	= partial_clause_prev[5][138] & 1'b1;
			partial_clause[5][139] 	= partial_clause_prev[5][139] & 1'b1;
			partial_clause[5][140] 	= partial_clause_prev[5][140] & 1'b1;
			partial_clause[5][141] 	= partial_clause_prev[5][141] & x[8];
			partial_clause[5][142] 	= partial_clause_prev[5][142] & 1'b1;
			partial_clause[5][143] 	= partial_clause_prev[5][143] & 1'b1;
			partial_clause[5][144] 	= partial_clause_prev[5][144] & 1'b1;
			partial_clause[5][145] 	= partial_clause_prev[5][145] & 1'b1;
			partial_clause[5][146] 	= partial_clause_prev[5][146] & x[11] & x[38];
			partial_clause[5][147] 	= partial_clause_prev[5][147] & 1'b1;
			partial_clause[5][148] 	= partial_clause_prev[5][148] & 1'b1;
			partial_clause[5][149] 	= partial_clause_prev[5][149] & 1'b1;
			partial_clause[5][150] 	= partial_clause_prev[5][150] & 1'b1;
			partial_clause[5][151] 	= partial_clause_prev[5][151] & x[16];
			partial_clause[5][152] 	= partial_clause_prev[5][152] & ~x[63];
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & 1'b1;
			partial_clause[5][155] 	= partial_clause_prev[5][155] & 1'b1;
			partial_clause[5][156] 	= partial_clause_prev[5][156] & 1'b1;
			partial_clause[5][157] 	= partial_clause_prev[5][157] & ~x[35];
			partial_clause[5][158] 	= partial_clause_prev[5][158] & x[41];
			partial_clause[5][159] 	= partial_clause_prev[5][159] & x[11];
			partial_clause[5][160] 	= partial_clause_prev[5][160] & 1'b1;
			partial_clause[5][161] 	= partial_clause_prev[5][161] & 1'b1;
			partial_clause[5][162] 	= partial_clause_prev[5][162] & x[8];
			partial_clause[5][163] 	= partial_clause_prev[5][163] & 1'b1;
			partial_clause[5][164] 	= partial_clause_prev[5][164] & ~x[62];
			partial_clause[5][165] 	= partial_clause_prev[5][165] & 1'b1;
			partial_clause[5][166] 	= partial_clause_prev[5][166] & 1'b1;
			partial_clause[5][167] 	= partial_clause_prev[5][167] & 1'b1;
			partial_clause[5][168] 	= partial_clause_prev[5][168] & 1'b1;
			partial_clause[5][169] 	= partial_clause_prev[5][169] & x[14] & ~x[34] & ~x[62];
			partial_clause[5][170] 	= partial_clause_prev[5][170] & 1'b1;
			partial_clause[5][171] 	= partial_clause_prev[5][171] & 1'b1;
			partial_clause[5][172] 	= partial_clause_prev[5][172] & 1'b1;
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & 1'b1;
			partial_clause[5][175] 	= partial_clause_prev[5][175] & 1'b1;
			partial_clause[5][176] 	= partial_clause_prev[5][176] & 1'b1;
			partial_clause[5][177] 	= partial_clause_prev[5][177] & ~x[6];
			partial_clause[5][178] 	= partial_clause_prev[5][178] & 1'b1;
			partial_clause[5][179] 	= partial_clause_prev[5][179] & 1'b1;
			partial_clause[5][180] 	= partial_clause_prev[5][180] & 1'b1;
			partial_clause[5][181] 	= partial_clause_prev[5][181] & 1'b1;
			partial_clause[5][182] 	= partial_clause_prev[5][182] & 1'b1;
			partial_clause[5][183] 	= partial_clause_prev[5][183] & x[14];
			partial_clause[5][184] 	= partial_clause_prev[5][184] & 1'b1;
			partial_clause[5][185] 	= partial_clause_prev[5][185] & 1'b1;
			partial_clause[5][186] 	= partial_clause_prev[5][186] & 1'b1;
			partial_clause[5][187] 	= partial_clause_prev[5][187] & 1'b1;
			partial_clause[5][188] 	= partial_clause_prev[5][188] & 1'b1;
			partial_clause[5][189] 	= partial_clause_prev[5][189] & ~x[63];
			partial_clause[5][190] 	= partial_clause_prev[5][190] & 1'b1;
			partial_clause[5][191] 	= partial_clause_prev[5][191] & 1'b1;
			partial_clause[5][192] 	= partial_clause_prev[5][192] & 1'b1;
			partial_clause[5][193] 	= partial_clause_prev[5][193] & 1'b1;
			partial_clause[5][194] 	= partial_clause_prev[5][194] & 1'b1;
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & 1'b1;
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & 1'b1;
			partial_clause[5][199] 	= partial_clause_prev[5][199] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & x[9];
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & ~x[32];
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & x[39];
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & x[9] & x[37];
			partial_clause[6][47] 	= partial_clause_prev[6][47] & x[12];
			partial_clause[6][48] 	= partial_clause_prev[6][48] & x[40];
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & x[19];
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & ~x[17];
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			partial_clause[6][100] 	= partial_clause_prev[6][100] & 1'b1;
			partial_clause[6][101] 	= partial_clause_prev[6][101] & 1'b1;
			partial_clause[6][102] 	= partial_clause_prev[6][102] & 1'b1;
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & 1'b1;
			partial_clause[6][105] 	= partial_clause_prev[6][105] & 1'b1;
			partial_clause[6][106] 	= partial_clause_prev[6][106] & 1'b1;
			partial_clause[6][107] 	= partial_clause_prev[6][107] & 1'b1;
			partial_clause[6][108] 	= partial_clause_prev[6][108] & 1'b1;
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & 1'b1;
			partial_clause[6][111] 	= partial_clause_prev[6][111] & ~x[63];
			partial_clause[6][112] 	= partial_clause_prev[6][112] & ~x[20];
			partial_clause[6][113] 	= partial_clause_prev[6][113] & 1'b1;
			partial_clause[6][114] 	= partial_clause_prev[6][114] & 1'b1;
			partial_clause[6][115] 	= partial_clause_prev[6][115] & 1'b1;
			partial_clause[6][116] 	= partial_clause_prev[6][116] & 1'b1;
			partial_clause[6][117] 	= partial_clause_prev[6][117] & 1'b1;
			partial_clause[6][118] 	= partial_clause_prev[6][118] & 1'b1;
			partial_clause[6][119] 	= partial_clause_prev[6][119] & 1'b1;
			partial_clause[6][120] 	= partial_clause_prev[6][120] & 1'b1;
			partial_clause[6][121] 	= partial_clause_prev[6][121] & 1'b1;
			partial_clause[6][122] 	= partial_clause_prev[6][122] & 1'b1;
			partial_clause[6][123] 	= partial_clause_prev[6][123] & ~x[38];
			partial_clause[6][124] 	= partial_clause_prev[6][124] & 1'b1;
			partial_clause[6][125] 	= partial_clause_prev[6][125] & 1'b1;
			partial_clause[6][126] 	= partial_clause_prev[6][126] & 1'b1;
			partial_clause[6][127] 	= partial_clause_prev[6][127] & 1'b1;
			partial_clause[6][128] 	= partial_clause_prev[6][128] & 1'b1;
			partial_clause[6][129] 	= partial_clause_prev[6][129] & 1'b1;
			partial_clause[6][130] 	= partial_clause_prev[6][130] & 1'b1;
			partial_clause[6][131] 	= partial_clause_prev[6][131] & 1'b1;
			partial_clause[6][132] 	= partial_clause_prev[6][132] & 1'b1;
			partial_clause[6][133] 	= partial_clause_prev[6][133] & 1'b1;
			partial_clause[6][134] 	= partial_clause_prev[6][134] & 1'b1;
			partial_clause[6][135] 	= partial_clause_prev[6][135] & 1'b1;
			partial_clause[6][136] 	= partial_clause_prev[6][136] & 1'b1;
			partial_clause[6][137] 	= partial_clause_prev[6][137] & 1'b1;
			partial_clause[6][138] 	= partial_clause_prev[6][138] & 1'b1;
			partial_clause[6][139] 	= partial_clause_prev[6][139] & 1'b1;
			partial_clause[6][140] 	= partial_clause_prev[6][140] & 1'b1;
			partial_clause[6][141] 	= partial_clause_prev[6][141] & 1'b1;
			partial_clause[6][142] 	= partial_clause_prev[6][142] & 1'b1;
			partial_clause[6][143] 	= partial_clause_prev[6][143] & 1'b1;
			partial_clause[6][144] 	= partial_clause_prev[6][144] & 1'b1;
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & 1'b1;
			partial_clause[6][147] 	= partial_clause_prev[6][147] & 1'b1;
			partial_clause[6][148] 	= partial_clause_prev[6][148] & 1'b1;
			partial_clause[6][149] 	= partial_clause_prev[6][149] & 1'b1;
			partial_clause[6][150] 	= partial_clause_prev[6][150] & 1'b1;
			partial_clause[6][151] 	= partial_clause_prev[6][151] & 1'b1;
			partial_clause[6][152] 	= partial_clause_prev[6][152] & 1'b1;
			partial_clause[6][153] 	= partial_clause_prev[6][153] & ~x[15];
			partial_clause[6][154] 	= partial_clause_prev[6][154] & 1'b1;
			partial_clause[6][155] 	= partial_clause_prev[6][155] & 1'b1;
			partial_clause[6][156] 	= partial_clause_prev[6][156] & 1'b1;
			partial_clause[6][157] 	= partial_clause_prev[6][157] & 1'b1;
			partial_clause[6][158] 	= partial_clause_prev[6][158] & ~x[7];
			partial_clause[6][159] 	= partial_clause_prev[6][159] & ~x[38];
			partial_clause[6][160] 	= partial_clause_prev[6][160] & ~x[6] & ~x[11];
			partial_clause[6][161] 	= partial_clause_prev[6][161] & 1'b1;
			partial_clause[6][162] 	= partial_clause_prev[6][162] & 1'b1;
			partial_clause[6][163] 	= partial_clause_prev[6][163] & 1'b1;
			partial_clause[6][164] 	= partial_clause_prev[6][164] & 1'b1;
			partial_clause[6][165] 	= partial_clause_prev[6][165] & 1'b1;
			partial_clause[6][166] 	= partial_clause_prev[6][166] & 1'b1;
			partial_clause[6][167] 	= partial_clause_prev[6][167] & 1'b1;
			partial_clause[6][168] 	= partial_clause_prev[6][168] & 1'b1;
			partial_clause[6][169] 	= partial_clause_prev[6][169] & ~x[6] & ~x[8] & ~x[9] & ~x[10];
			partial_clause[6][170] 	= partial_clause_prev[6][170] & 1'b1;
			partial_clause[6][171] 	= partial_clause_prev[6][171] & 1'b1;
			partial_clause[6][172] 	= partial_clause_prev[6][172] & ~x[7] & ~x[11] & ~x[37];
			partial_clause[6][173] 	= partial_clause_prev[6][173] & 1'b1;
			partial_clause[6][174] 	= partial_clause_prev[6][174] & 1'b1;
			partial_clause[6][175] 	= partial_clause_prev[6][175] & 1'b1;
			partial_clause[6][176] 	= partial_clause_prev[6][176] & 1'b1;
			partial_clause[6][177] 	= partial_clause_prev[6][177] & 1'b1;
			partial_clause[6][178] 	= partial_clause_prev[6][178] & 1'b1;
			partial_clause[6][179] 	= partial_clause_prev[6][179] & 1'b1;
			partial_clause[6][180] 	= partial_clause_prev[6][180] & 1'b1;
			partial_clause[6][181] 	= partial_clause_prev[6][181] & 1'b1;
			partial_clause[6][182] 	= partial_clause_prev[6][182] & 1'b1;
			partial_clause[6][183] 	= partial_clause_prev[6][183] & ~x[9] & ~x[11];
			partial_clause[6][184] 	= partial_clause_prev[6][184] & 1'b1;
			partial_clause[6][185] 	= partial_clause_prev[6][185] & ~x[37] & ~x[39] & ~x[63];
			partial_clause[6][186] 	= partial_clause_prev[6][186] & 1'b1;
			partial_clause[6][187] 	= partial_clause_prev[6][187] & 1'b1;
			partial_clause[6][188] 	= partial_clause_prev[6][188] & 1'b1;
			partial_clause[6][189] 	= partial_clause_prev[6][189] & 1'b1;
			partial_clause[6][190] 	= partial_clause_prev[6][190] & 1'b1;
			partial_clause[6][191] 	= partial_clause_prev[6][191] & 1'b1;
			partial_clause[6][192] 	= partial_clause_prev[6][192] & 1'b1;
			partial_clause[6][193] 	= partial_clause_prev[6][193] & ~x[36] & ~x[37] & ~x[38] & ~x[39];
			partial_clause[6][194] 	= partial_clause_prev[6][194] & 1'b1;
			partial_clause[6][195] 	= partial_clause_prev[6][195] & 1'b1;
			partial_clause[6][196] 	= partial_clause_prev[6][196] & 1'b1;
			partial_clause[6][197] 	= partial_clause_prev[6][197] & ~x[9];
			partial_clause[6][198] 	= partial_clause_prev[6][198] & 1'b1;
			partial_clause[6][199] 	= partial_clause_prev[6][199] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & ~x[7];
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & ~x[12];
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & ~x[9] & ~x[63];
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & ~x[9];
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & ~x[40];
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & x[41];
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & ~x[13] & ~x[39];
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & x[42];
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & x[42];
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & x[16];
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & x[41];
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & ~x[38];
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & ~x[11];
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & x[42];
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & ~x[12];
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & ~x[11] & ~x[37];
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			partial_clause[7][100] 	= partial_clause_prev[7][100] & ~x[17];
			partial_clause[7][101] 	= partial_clause_prev[7][101] & ~x[19];
			partial_clause[7][102] 	= partial_clause_prev[7][102] & 1'b1;
			partial_clause[7][103] 	= partial_clause_prev[7][103] & 1'b1;
			partial_clause[7][104] 	= partial_clause_prev[7][104] & 1'b1;
			partial_clause[7][105] 	= partial_clause_prev[7][105] & 1'b1;
			partial_clause[7][106] 	= partial_clause_prev[7][106] & 1'b1;
			partial_clause[7][107] 	= partial_clause_prev[7][107] & x[62];
			partial_clause[7][108] 	= partial_clause_prev[7][108] & 1'b1;
			partial_clause[7][109] 	= partial_clause_prev[7][109] & 1'b1;
			partial_clause[7][110] 	= partial_clause_prev[7][110] & 1'b1;
			partial_clause[7][111] 	= partial_clause_prev[7][111] & 1'b1;
			partial_clause[7][112] 	= partial_clause_prev[7][112] & 1'b1;
			partial_clause[7][113] 	= partial_clause_prev[7][113] & 1'b1;
			partial_clause[7][114] 	= partial_clause_prev[7][114] & 1'b1;
			partial_clause[7][115] 	= partial_clause_prev[7][115] & 1'b1;
			partial_clause[7][116] 	= partial_clause_prev[7][116] & 1'b1;
			partial_clause[7][117] 	= partial_clause_prev[7][117] & 1'b1;
			partial_clause[7][118] 	= partial_clause_prev[7][118] & 1'b1;
			partial_clause[7][119] 	= partial_clause_prev[7][119] & 1'b1;
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & x[10];
			partial_clause[7][123] 	= partial_clause_prev[7][123] & 1'b1;
			partial_clause[7][124] 	= partial_clause_prev[7][124] & x[38];
			partial_clause[7][125] 	= partial_clause_prev[7][125] & 1'b1;
			partial_clause[7][126] 	= partial_clause_prev[7][126] & 1'b1;
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & 1'b1;
			partial_clause[7][129] 	= partial_clause_prev[7][129] & 1'b1;
			partial_clause[7][130] 	= partial_clause_prev[7][130] & 1'b1;
			partial_clause[7][131] 	= partial_clause_prev[7][131] & 1'b1;
			partial_clause[7][132] 	= partial_clause_prev[7][132] & 1'b1;
			partial_clause[7][133] 	= partial_clause_prev[7][133] & x[38];
			partial_clause[7][134] 	= partial_clause_prev[7][134] & 1'b1;
			partial_clause[7][135] 	= partial_clause_prev[7][135] & 1'b1;
			partial_clause[7][136] 	= partial_clause_prev[7][136] & x[11];
			partial_clause[7][137] 	= partial_clause_prev[7][137] & 1'b1;
			partial_clause[7][138] 	= partial_clause_prev[7][138] & x[8];
			partial_clause[7][139] 	= partial_clause_prev[7][139] & x[11];
			partial_clause[7][140] 	= partial_clause_prev[7][140] & 1'b1;
			partial_clause[7][141] 	= partial_clause_prev[7][141] & 1'b1;
			partial_clause[7][142] 	= partial_clause_prev[7][142] & 1'b1;
			partial_clause[7][143] 	= partial_clause_prev[7][143] & 1'b1;
			partial_clause[7][144] 	= partial_clause_prev[7][144] & 1'b1;
			partial_clause[7][145] 	= partial_clause_prev[7][145] & 1'b1;
			partial_clause[7][146] 	= partial_clause_prev[7][146] & ~x[18] & ~x[58];
			partial_clause[7][147] 	= partial_clause_prev[7][147] & 1'b1;
			partial_clause[7][148] 	= partial_clause_prev[7][148] & 1'b1;
			partial_clause[7][149] 	= partial_clause_prev[7][149] & 1'b1;
			partial_clause[7][150] 	= partial_clause_prev[7][150] & 1'b1;
			partial_clause[7][151] 	= partial_clause_prev[7][151] & 1'b1;
			partial_clause[7][152] 	= partial_clause_prev[7][152] & 1'b1;
			partial_clause[7][153] 	= partial_clause_prev[7][153] & 1'b1;
			partial_clause[7][154] 	= partial_clause_prev[7][154] & 1'b1;
			partial_clause[7][155] 	= partial_clause_prev[7][155] & 1'b1;
			partial_clause[7][156] 	= partial_clause_prev[7][156] & 1'b1;
			partial_clause[7][157] 	= partial_clause_prev[7][157] & 1'b1;
			partial_clause[7][158] 	= partial_clause_prev[7][158] & 1'b1;
			partial_clause[7][159] 	= partial_clause_prev[7][159] & 1'b1;
			partial_clause[7][160] 	= partial_clause_prev[7][160] & 1'b1;
			partial_clause[7][161] 	= partial_clause_prev[7][161] & 1'b1;
			partial_clause[7][162] 	= partial_clause_prev[7][162] & 1'b1;
			partial_clause[7][163] 	= partial_clause_prev[7][163] & x[10];
			partial_clause[7][164] 	= partial_clause_prev[7][164] & 1'b1;
			partial_clause[7][165] 	= partial_clause_prev[7][165] & 1'b1;
			partial_clause[7][166] 	= partial_clause_prev[7][166] & 1'b1;
			partial_clause[7][167] 	= partial_clause_prev[7][167] & 1'b1;
			partial_clause[7][168] 	= partial_clause_prev[7][168] & 1'b1;
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & 1'b1;
			partial_clause[7][171] 	= partial_clause_prev[7][171] & ~x[9];
			partial_clause[7][172] 	= partial_clause_prev[7][172] & ~x[6] & ~x[40];
			partial_clause[7][173] 	= partial_clause_prev[7][173] & x[10];
			partial_clause[7][174] 	= partial_clause_prev[7][174] & 1'b1;
			partial_clause[7][175] 	= partial_clause_prev[7][175] & 1'b1;
			partial_clause[7][176] 	= partial_clause_prev[7][176] & 1'b1;
			partial_clause[7][177] 	= partial_clause_prev[7][177] & 1'b1;
			partial_clause[7][178] 	= partial_clause_prev[7][178] & 1'b1;
			partial_clause[7][179] 	= partial_clause_prev[7][179] & ~x[41];
			partial_clause[7][180] 	= partial_clause_prev[7][180] & 1'b1;
			partial_clause[7][181] 	= partial_clause_prev[7][181] & 1'b1;
			partial_clause[7][182] 	= partial_clause_prev[7][182] & 1'b1;
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & 1'b1;
			partial_clause[7][185] 	= partial_clause_prev[7][185] & ~x[5] & ~x[8];
			partial_clause[7][186] 	= partial_clause_prev[7][186] & 1'b1;
			partial_clause[7][187] 	= partial_clause_prev[7][187] & 1'b1;
			partial_clause[7][188] 	= partial_clause_prev[7][188] & 1'b1;
			partial_clause[7][189] 	= partial_clause_prev[7][189] & 1'b1;
			partial_clause[7][190] 	= partial_clause_prev[7][190] & ~x[11];
			partial_clause[7][191] 	= partial_clause_prev[7][191] & 1'b1;
			partial_clause[7][192] 	= partial_clause_prev[7][192] & 1'b1;
			partial_clause[7][193] 	= partial_clause_prev[7][193] & 1'b1;
			partial_clause[7][194] 	= partial_clause_prev[7][194] & 1'b1;
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & ~x[58];
			partial_clause[7][197] 	= partial_clause_prev[7][197] & x[12];
			partial_clause[7][198] 	= partial_clause_prev[7][198] & 1'b1;
			partial_clause[7][199] 	= partial_clause_prev[7][199] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & x[39] & ~x[46];
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & ~x[8] & ~x[62];
			partial_clause[8][11] 	= partial_clause_prev[8][11] & ~x[20];
			partial_clause[8][12] 	= partial_clause_prev[8][12] & x[13] & x[40];
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & ~x[37];
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & ~x[8];
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & ~x[8] & ~x[37];
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & ~x[46];
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & ~x[46];
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & x[37];
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & x[39];
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & x[28];
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & ~x[37] & x[40];
			partial_clause[8][70] 	= partial_clause_prev[8][70] & x[37];
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & ~x[19] & ~x[36] & ~x[47];
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & x[13];
			partial_clause[8][82] 	= partial_clause_prev[8][82] & x[37];
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & ~x[36];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & x[1];
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & x[38];
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			partial_clause[8][100] 	= partial_clause_prev[8][100] & 1'b1;
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & 1'b1;
			partial_clause[8][103] 	= partial_clause_prev[8][103] & 1'b1;
			partial_clause[8][104] 	= partial_clause_prev[8][104] & 1'b1;
			partial_clause[8][105] 	= partial_clause_prev[8][105] & 1'b1;
			partial_clause[8][106] 	= partial_clause_prev[8][106] & x[7];
			partial_clause[8][107] 	= partial_clause_prev[8][107] & 1'b1;
			partial_clause[8][108] 	= partial_clause_prev[8][108] & x[4];
			partial_clause[8][109] 	= partial_clause_prev[8][109] & ~x[35] & ~x[36] & ~x[38];
			partial_clause[8][110] 	= partial_clause_prev[8][110] & 1'b1;
			partial_clause[8][111] 	= partial_clause_prev[8][111] & 1'b1;
			partial_clause[8][112] 	= partial_clause_prev[8][112] & 1'b1;
			partial_clause[8][113] 	= partial_clause_prev[8][113] & 1'b1;
			partial_clause[8][114] 	= partial_clause_prev[8][114] & 1'b1;
			partial_clause[8][115] 	= partial_clause_prev[8][115] & 1'b1;
			partial_clause[8][116] 	= partial_clause_prev[8][116] & 1'b1;
			partial_clause[8][117] 	= partial_clause_prev[8][117] & 1'b1;
			partial_clause[8][118] 	= partial_clause_prev[8][118] & ~x[10] & ~x[12] & ~x[13];
			partial_clause[8][119] 	= partial_clause_prev[8][119] & ~x[35];
			partial_clause[8][120] 	= partial_clause_prev[8][120] & 1'b1;
			partial_clause[8][121] 	= partial_clause_prev[8][121] & 1'b1;
			partial_clause[8][122] 	= partial_clause_prev[8][122] & 1'b1;
			partial_clause[8][123] 	= partial_clause_prev[8][123] & 1'b1;
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & 1'b1;
			partial_clause[8][126] 	= partial_clause_prev[8][126] & 1'b1;
			partial_clause[8][127] 	= partial_clause_prev[8][127] & 1'b1;
			partial_clause[8][128] 	= partial_clause_prev[8][128] & x[18];
			partial_clause[8][129] 	= partial_clause_prev[8][129] & ~x[8] & ~x[13];
			partial_clause[8][130] 	= partial_clause_prev[8][130] & ~x[39] & ~x[41];
			partial_clause[8][131] 	= partial_clause_prev[8][131] & 1'b1;
			partial_clause[8][132] 	= partial_clause_prev[8][132] & 1'b1;
			partial_clause[8][133] 	= partial_clause_prev[8][133] & 1'b1;
			partial_clause[8][134] 	= partial_clause_prev[8][134] & 1'b1;
			partial_clause[8][135] 	= partial_clause_prev[8][135] & 1'b1;
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & 1'b1;
			partial_clause[8][138] 	= partial_clause_prev[8][138] & 1'b1;
			partial_clause[8][139] 	= partial_clause_prev[8][139] & 1'b1;
			partial_clause[8][140] 	= partial_clause_prev[8][140] & 1'b1;
			partial_clause[8][141] 	= partial_clause_prev[8][141] & 1'b1;
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & ~x[12] & ~x[13];
			partial_clause[8][144] 	= partial_clause_prev[8][144] & x[22];
			partial_clause[8][145] 	= partial_clause_prev[8][145] & 1'b1;
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & 1'b1;
			partial_clause[8][148] 	= partial_clause_prev[8][148] & x[19];
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & 1'b1;
			partial_clause[8][151] 	= partial_clause_prev[8][151] & 1'b1;
			partial_clause[8][152] 	= partial_clause_prev[8][152] & ~x[34];
			partial_clause[8][153] 	= partial_clause_prev[8][153] & 1'b1;
			partial_clause[8][154] 	= partial_clause_prev[8][154] & 1'b1;
			partial_clause[8][155] 	= partial_clause_prev[8][155] & ~x[2] & ~x[7] & ~x[8] & ~x[38] & ~x[40];
			partial_clause[8][156] 	= partial_clause_prev[8][156] & 1'b1;
			partial_clause[8][157] 	= partial_clause_prev[8][157] & 1'b1;
			partial_clause[8][158] 	= partial_clause_prev[8][158] & 1'b1;
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & 1'b1;
			partial_clause[8][161] 	= partial_clause_prev[8][161] & 1'b1;
			partial_clause[8][162] 	= partial_clause_prev[8][162] & 1'b1;
			partial_clause[8][163] 	= partial_clause_prev[8][163] & 1'b1;
			partial_clause[8][164] 	= partial_clause_prev[8][164] & 1'b1;
			partial_clause[8][165] 	= partial_clause_prev[8][165] & 1'b1;
			partial_clause[8][166] 	= partial_clause_prev[8][166] & ~x[7] & ~x[39];
			partial_clause[8][167] 	= partial_clause_prev[8][167] & x[17];
			partial_clause[8][168] 	= partial_clause_prev[8][168] & 1'b1;
			partial_clause[8][169] 	= partial_clause_prev[8][169] & 1'b1;
			partial_clause[8][170] 	= partial_clause_prev[8][170] & 1'b1;
			partial_clause[8][171] 	= partial_clause_prev[8][171] & 1'b1;
			partial_clause[8][172] 	= partial_clause_prev[8][172] & 1'b1;
			partial_clause[8][173] 	= partial_clause_prev[8][173] & 1'b1;
			partial_clause[8][174] 	= partial_clause_prev[8][174] & 1'b1;
			partial_clause[8][175] 	= partial_clause_prev[8][175] & 1'b1;
			partial_clause[8][176] 	= partial_clause_prev[8][176] & 1'b1;
			partial_clause[8][177] 	= partial_clause_prev[8][177] & x[36];
			partial_clause[8][178] 	= partial_clause_prev[8][178] & 1'b1;
			partial_clause[8][179] 	= partial_clause_prev[8][179] & 1'b1;
			partial_clause[8][180] 	= partial_clause_prev[8][180] & 1'b1;
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & 1'b1;
			partial_clause[8][183] 	= partial_clause_prev[8][183] & 1'b1;
			partial_clause[8][184] 	= partial_clause_prev[8][184] & 1'b1;
			partial_clause[8][185] 	= partial_clause_prev[8][185] & 1'b1;
			partial_clause[8][186] 	= partial_clause_prev[8][186] & 1'b1;
			partial_clause[8][187] 	= partial_clause_prev[8][187] & 1'b1;
			partial_clause[8][188] 	= partial_clause_prev[8][188] & ~x[16];
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & ~x[63];
			partial_clause[8][191] 	= partial_clause_prev[8][191] & x[54];
			partial_clause[8][192] 	= partial_clause_prev[8][192] & ~x[44];
			partial_clause[8][193] 	= partial_clause_prev[8][193] & 1'b1;
			partial_clause[8][194] 	= partial_clause_prev[8][194] & 1'b1;
			partial_clause[8][195] 	= partial_clause_prev[8][195] & 1'b1;
			partial_clause[8][196] 	= partial_clause_prev[8][196] & 1'b1;
			partial_clause[8][197] 	= partial_clause_prev[8][197] & 1'b1;
			partial_clause[8][198] 	= partial_clause_prev[8][198] & 1'b1;
			partial_clause[8][199] 	= partial_clause_prev[8][199] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & ~x[51];
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & x[16] & ~x[22] & ~x[47];
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & x[16];
			partial_clause[9][35] 	= partial_clause_prev[9][35] & 1'b1;
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & ~x[41];
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & ~x[47];
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & ~x[19];
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & ~x[47];
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & ~x[47];
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & ~x[20];
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & ~x[20];
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & ~x[21];
			partial_clause[9][100] 	= partial_clause_prev[9][100] & 1'b1;
			partial_clause[9][101] 	= partial_clause_prev[9][101] & 1'b1;
			partial_clause[9][102] 	= partial_clause_prev[9][102] & x[13];
			partial_clause[9][103] 	= partial_clause_prev[9][103] & 1'b1;
			partial_clause[9][104] 	= partial_clause_prev[9][104] & 1'b1;
			partial_clause[9][105] 	= partial_clause_prev[9][105] & x[21];
			partial_clause[9][106] 	= partial_clause_prev[9][106] & 1'b1;
			partial_clause[9][107] 	= partial_clause_prev[9][107] & 1'b1;
			partial_clause[9][108] 	= partial_clause_prev[9][108] & 1'b1;
			partial_clause[9][109] 	= partial_clause_prev[9][109] & 1'b1;
			partial_clause[9][110] 	= partial_clause_prev[9][110] & 1'b1;
			partial_clause[9][111] 	= partial_clause_prev[9][111] & 1'b1;
			partial_clause[9][112] 	= partial_clause_prev[9][112] & 1'b1;
			partial_clause[9][113] 	= partial_clause_prev[9][113] & 1'b1;
			partial_clause[9][114] 	= partial_clause_prev[9][114] & 1'b1;
			partial_clause[9][115] 	= partial_clause_prev[9][115] & 1'b1;
			partial_clause[9][116] 	= partial_clause_prev[9][116] & ~x[40];
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & 1'b1;
			partial_clause[9][119] 	= partial_clause_prev[9][119] & 1'b1;
			partial_clause[9][120] 	= partial_clause_prev[9][120] & 1'b1;
			partial_clause[9][121] 	= partial_clause_prev[9][121] & 1'b1;
			partial_clause[9][122] 	= partial_clause_prev[9][122] & 1'b1;
			partial_clause[9][123] 	= partial_clause_prev[9][123] & 1'b1;
			partial_clause[9][124] 	= partial_clause_prev[9][124] & 1'b1;
			partial_clause[9][125] 	= partial_clause_prev[9][125] & 1'b1;
			partial_clause[9][126] 	= partial_clause_prev[9][126] & 1'b1;
			partial_clause[9][127] 	= partial_clause_prev[9][127] & 1'b1;
			partial_clause[9][128] 	= partial_clause_prev[9][128] & 1'b1;
			partial_clause[9][129] 	= partial_clause_prev[9][129] & 1'b1;
			partial_clause[9][130] 	= partial_clause_prev[9][130] & 1'b1;
			partial_clause[9][131] 	= partial_clause_prev[9][131] & 1'b1;
			partial_clause[9][132] 	= partial_clause_prev[9][132] & 1'b1;
			partial_clause[9][133] 	= partial_clause_prev[9][133] & x[39];
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & 1'b1;
			partial_clause[9][138] 	= partial_clause_prev[9][138] & 1'b1;
			partial_clause[9][139] 	= partial_clause_prev[9][139] & 1'b1;
			partial_clause[9][140] 	= partial_clause_prev[9][140] & 1'b1;
			partial_clause[9][141] 	= partial_clause_prev[9][141] & 1'b1;
			partial_clause[9][142] 	= partial_clause_prev[9][142] & 1'b1;
			partial_clause[9][143] 	= partial_clause_prev[9][143] & x[21];
			partial_clause[9][144] 	= partial_clause_prev[9][144] & 1'b1;
			partial_clause[9][145] 	= partial_clause_prev[9][145] & 1'b1;
			partial_clause[9][146] 	= partial_clause_prev[9][146] & 1'b1;
			partial_clause[9][147] 	= partial_clause_prev[9][147] & 1'b1;
			partial_clause[9][148] 	= partial_clause_prev[9][148] & ~x[8] & ~x[34];
			partial_clause[9][149] 	= partial_clause_prev[9][149] & 1'b1;
			partial_clause[9][150] 	= partial_clause_prev[9][150] & x[50];
			partial_clause[9][151] 	= partial_clause_prev[9][151] & 1'b1;
			partial_clause[9][152] 	= partial_clause_prev[9][152] & 1'b1;
			partial_clause[9][153] 	= partial_clause_prev[9][153] & 1'b1;
			partial_clause[9][154] 	= partial_clause_prev[9][154] & 1'b1;
			partial_clause[9][155] 	= partial_clause_prev[9][155] & 1'b1;
			partial_clause[9][156] 	= partial_clause_prev[9][156] & 1'b1;
			partial_clause[9][157] 	= partial_clause_prev[9][157] & 1'b1;
			partial_clause[9][158] 	= partial_clause_prev[9][158] & 1'b1;
			partial_clause[9][159] 	= partial_clause_prev[9][159] & 1'b1;
			partial_clause[9][160] 	= partial_clause_prev[9][160] & 1'b1;
			partial_clause[9][161] 	= partial_clause_prev[9][161] & x[49];
			partial_clause[9][162] 	= partial_clause_prev[9][162] & 1'b1;
			partial_clause[9][163] 	= partial_clause_prev[9][163] & 1'b1;
			partial_clause[9][164] 	= partial_clause_prev[9][164] & 1'b1;
			partial_clause[9][165] 	= partial_clause_prev[9][165] & 1'b1;
			partial_clause[9][166] 	= partial_clause_prev[9][166] & 1'b1;
			partial_clause[9][167] 	= partial_clause_prev[9][167] & ~x[10] & ~x[36] & ~x[63];
			partial_clause[9][168] 	= partial_clause_prev[9][168] & 1'b1;
			partial_clause[9][169] 	= partial_clause_prev[9][169] & 1'b1;
			partial_clause[9][170] 	= partial_clause_prev[9][170] & ~x[18];
			partial_clause[9][171] 	= partial_clause_prev[9][171] & 1'b1;
			partial_clause[9][172] 	= partial_clause_prev[9][172] & ~x[6];
			partial_clause[9][173] 	= partial_clause_prev[9][173] & 1'b1;
			partial_clause[9][174] 	= partial_clause_prev[9][174] & 1'b1;
			partial_clause[9][175] 	= partial_clause_prev[9][175] & 1'b1;
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & 1'b1;
			partial_clause[9][178] 	= partial_clause_prev[9][178] & 1'b1;
			partial_clause[9][179] 	= partial_clause_prev[9][179] & 1'b1;
			partial_clause[9][180] 	= partial_clause_prev[9][180] & 1'b1;
			partial_clause[9][181] 	= partial_clause_prev[9][181] & 1'b1;
			partial_clause[9][182] 	= partial_clause_prev[9][182] & 1'b1;
			partial_clause[9][183] 	= partial_clause_prev[9][183] & 1'b1;
			partial_clause[9][184] 	= partial_clause_prev[9][184] & 1'b1;
			partial_clause[9][185] 	= partial_clause_prev[9][185] & 1'b1;
			partial_clause[9][186] 	= partial_clause_prev[9][186] & 1'b1;
			partial_clause[9][187] 	= partial_clause_prev[9][187] & 1'b1;
			partial_clause[9][188] 	= partial_clause_prev[9][188] & 1'b1;
			partial_clause[9][189] 	= partial_clause_prev[9][189] & 1'b1;
			partial_clause[9][190] 	= partial_clause_prev[9][190] & 1'b1;
			partial_clause[9][191] 	= partial_clause_prev[9][191] & 1'b1;
			partial_clause[9][192] 	= partial_clause_prev[9][192] & 1'b1;
			partial_clause[9][193] 	= partial_clause_prev[9][193] & 1'b1;
			partial_clause[9][194] 	= partial_clause_prev[9][194] & 1'b1;
			partial_clause[9][195] 	= partial_clause_prev[9][195] & 1'b1;
			partial_clause[9][196] 	= partial_clause_prev[9][196] & ~x[7] & ~x[8];
			partial_clause[9][197] 	= partial_clause_prev[9][197] & 1'b1;
			partial_clause[9][198] 	= partial_clause_prev[9][198] & 1'b1;
			partial_clause[9][199] 	= partial_clause_prev[9][199] & 1'b1;
		end
	end
endmodule


module HCB_8 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & ~x[5];
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & x[57];
			partial_clause[0][3] 	= partial_clause_prev[0][3] & x[57];
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & ~x[7];
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & x[8] & ~x[39];
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & ~x[34];
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & ~x[40];
			partial_clause[0][16] 	= partial_clause_prev[0][16] & x[0] & ~x[3] & ~x[40];
			partial_clause[0][17] 	= partial_clause_prev[0][17] & x[28];
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & x[0];
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & x[2] & ~x[25];
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & x[28];
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & x[56];
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & x[0];
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & x[1] & ~x[26];
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & ~x[7];
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & x[59];
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & ~x[8] & ~x[35];
			partial_clause[0][65] 	= partial_clause_prev[0][65] & ~x[6];
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & x[30] & ~x[54];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & x[2] & ~x[55];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & ~x[32];
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & x[20];
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & x[30];
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & x[27];
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			partial_clause[0][100] 	= partial_clause_prev[0][100] & 1'b1;
			partial_clause[0][101] 	= partial_clause_prev[0][101] & 1'b1;
			partial_clause[0][102] 	= partial_clause_prev[0][102] & 1'b1;
			partial_clause[0][103] 	= partial_clause_prev[0][103] & 1'b1;
			partial_clause[0][104] 	= partial_clause_prev[0][104] & 1'b1;
			partial_clause[0][105] 	= partial_clause_prev[0][105] & ~x[28] & ~x[58];
			partial_clause[0][106] 	= partial_clause_prev[0][106] & 1'b1;
			partial_clause[0][107] 	= partial_clause_prev[0][107] & 1'b1;
			partial_clause[0][108] 	= partial_clause_prev[0][108] & ~x[57];
			partial_clause[0][109] 	= partial_clause_prev[0][109] & 1'b1;
			partial_clause[0][110] 	= partial_clause_prev[0][110] & 1'b1;
			partial_clause[0][111] 	= partial_clause_prev[0][111] & 1'b1;
			partial_clause[0][112] 	= partial_clause_prev[0][112] & 1'b1;
			partial_clause[0][113] 	= partial_clause_prev[0][113] & 1'b1;
			partial_clause[0][114] 	= partial_clause_prev[0][114] & 1'b1;
			partial_clause[0][115] 	= partial_clause_prev[0][115] & 1'b1;
			partial_clause[0][116] 	= partial_clause_prev[0][116] & x[35];
			partial_clause[0][117] 	= partial_clause_prev[0][117] & x[63];
			partial_clause[0][118] 	= partial_clause_prev[0][118] & 1'b1;
			partial_clause[0][119] 	= partial_clause_prev[0][119] & 1'b1;
			partial_clause[0][120] 	= partial_clause_prev[0][120] & 1'b1;
			partial_clause[0][121] 	= partial_clause_prev[0][121] & 1'b1;
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & 1'b1;
			partial_clause[0][124] 	= partial_clause_prev[0][124] & 1'b1;
			partial_clause[0][125] 	= partial_clause_prev[0][125] & 1'b1;
			partial_clause[0][126] 	= partial_clause_prev[0][126] & ~x[3];
			partial_clause[0][127] 	= partial_clause_prev[0][127] & 1'b1;
			partial_clause[0][128] 	= partial_clause_prev[0][128] & ~x[30];
			partial_clause[0][129] 	= partial_clause_prev[0][129] & 1'b1;
			partial_clause[0][130] 	= partial_clause_prev[0][130] & ~x[31];
			partial_clause[0][131] 	= partial_clause_prev[0][131] & 1'b1;
			partial_clause[0][132] 	= partial_clause_prev[0][132] & 1'b1;
			partial_clause[0][133] 	= partial_clause_prev[0][133] & 1'b1;
			partial_clause[0][134] 	= partial_clause_prev[0][134] & 1'b1;
			partial_clause[0][135] 	= partial_clause_prev[0][135] & 1'b1;
			partial_clause[0][136] 	= partial_clause_prev[0][136] & 1'b1;
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & ~x[1] & ~x[26];
			partial_clause[0][139] 	= partial_clause_prev[0][139] & 1'b1;
			partial_clause[0][140] 	= partial_clause_prev[0][140] & 1'b1;
			partial_clause[0][141] 	= partial_clause_prev[0][141] & 1'b1;
			partial_clause[0][142] 	= partial_clause_prev[0][142] & ~x[2];
			partial_clause[0][143] 	= partial_clause_prev[0][143] & 1'b1;
			partial_clause[0][144] 	= partial_clause_prev[0][144] & 1'b1;
			partial_clause[0][145] 	= partial_clause_prev[0][145] & 1'b1;
			partial_clause[0][146] 	= partial_clause_prev[0][146] & 1'b1;
			partial_clause[0][147] 	= partial_clause_prev[0][147] & x[9];
			partial_clause[0][148] 	= partial_clause_prev[0][148] & 1'b1;
			partial_clause[0][149] 	= partial_clause_prev[0][149] & x[63];
			partial_clause[0][150] 	= partial_clause_prev[0][150] & 1'b1;
			partial_clause[0][151] 	= partial_clause_prev[0][151] & 1'b1;
			partial_clause[0][152] 	= partial_clause_prev[0][152] & 1'b1;
			partial_clause[0][153] 	= partial_clause_prev[0][153] & ~x[28] & ~x[29] & ~x[30];
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & 1'b1;
			partial_clause[0][156] 	= partial_clause_prev[0][156] & 1'b1;
			partial_clause[0][157] 	= partial_clause_prev[0][157] & 1'b1;
			partial_clause[0][158] 	= partial_clause_prev[0][158] & 1'b1;
			partial_clause[0][159] 	= partial_clause_prev[0][159] & 1'b1;
			partial_clause[0][160] 	= partial_clause_prev[0][160] & x[23];
			partial_clause[0][161] 	= partial_clause_prev[0][161] & x[63];
			partial_clause[0][162] 	= partial_clause_prev[0][162] & ~x[32];
			partial_clause[0][163] 	= partial_clause_prev[0][163] & 1'b1;
			partial_clause[0][164] 	= partial_clause_prev[0][164] & 1'b1;
			partial_clause[0][165] 	= partial_clause_prev[0][165] & ~x[59];
			partial_clause[0][166] 	= partial_clause_prev[0][166] & 1'b1;
			partial_clause[0][167] 	= partial_clause_prev[0][167] & x[38];
			partial_clause[0][168] 	= partial_clause_prev[0][168] & 1'b1;
			partial_clause[0][169] 	= partial_clause_prev[0][169] & 1'b1;
			partial_clause[0][170] 	= partial_clause_prev[0][170] & 1'b1;
			partial_clause[0][171] 	= partial_clause_prev[0][171] & 1'b1;
			partial_clause[0][172] 	= partial_clause_prev[0][172] & 1'b1;
			partial_clause[0][173] 	= partial_clause_prev[0][173] & 1'b1;
			partial_clause[0][174] 	= partial_clause_prev[0][174] & 1'b1;
			partial_clause[0][175] 	= partial_clause_prev[0][175] & 1'b1;
			partial_clause[0][176] 	= partial_clause_prev[0][176] & 1'b1;
			partial_clause[0][177] 	= partial_clause_prev[0][177] & 1'b1;
			partial_clause[0][178] 	= partial_clause_prev[0][178] & 1'b1;
			partial_clause[0][179] 	= partial_clause_prev[0][179] & 1'b1;
			partial_clause[0][180] 	= partial_clause_prev[0][180] & 1'b1;
			partial_clause[0][181] 	= partial_clause_prev[0][181] & 1'b1;
			partial_clause[0][182] 	= partial_clause_prev[0][182] & 1'b1;
			partial_clause[0][183] 	= partial_clause_prev[0][183] & 1'b1;
			partial_clause[0][184] 	= partial_clause_prev[0][184] & ~x[2];
			partial_clause[0][185] 	= partial_clause_prev[0][185] & 1'b1;
			partial_clause[0][186] 	= partial_clause_prev[0][186] & 1'b1;
			partial_clause[0][187] 	= partial_clause_prev[0][187] & 1'b1;
			partial_clause[0][188] 	= partial_clause_prev[0][188] & 1'b1;
			partial_clause[0][189] 	= partial_clause_prev[0][189] & ~x[21];
			partial_clause[0][190] 	= partial_clause_prev[0][190] & 1'b1;
			partial_clause[0][191] 	= partial_clause_prev[0][191] & 1'b1;
			partial_clause[0][192] 	= partial_clause_prev[0][192] & 1'b1;
			partial_clause[0][193] 	= partial_clause_prev[0][193] & 1'b1;
			partial_clause[0][194] 	= partial_clause_prev[0][194] & 1'b1;
			partial_clause[0][195] 	= partial_clause_prev[0][195] & 1'b1;
			partial_clause[0][196] 	= partial_clause_prev[0][196] & ~x[0] & ~x[25] & ~x[53];
			partial_clause[0][197] 	= partial_clause_prev[0][197] & 1'b1;
			partial_clause[0][198] 	= partial_clause_prev[0][198] & 1'b1;
			partial_clause[0][199] 	= partial_clause_prev[0][199] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[7];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & x[6] & x[34];
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & ~x[10] & ~x[35];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & x[35];
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & ~x[2] & x[7] & x[35];
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & ~x[30];
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & x[34];
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & ~x[8];
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & x[31];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & ~x[34];
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & ~x[41];
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & x[48];
			partial_clause[1][74] 	= partial_clause_prev[1][74] & x[33];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & ~x[37] & ~x[63];
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & ~x[9] & x[60];
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & ~x[31] & ~x[58];
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & ~x[9];
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & x[47];
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & ~x[36];
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			partial_clause[1][100] 	= partial_clause_prev[1][100] & 1'b1;
			partial_clause[1][101] 	= partial_clause_prev[1][101] & 1'b1;
			partial_clause[1][102] 	= partial_clause_prev[1][102] & 1'b1;
			partial_clause[1][103] 	= partial_clause_prev[1][103] & 1'b1;
			partial_clause[1][104] 	= partial_clause_prev[1][104] & 1'b1;
			partial_clause[1][105] 	= partial_clause_prev[1][105] & 1'b1;
			partial_clause[1][106] 	= partial_clause_prev[1][106] & 1'b1;
			partial_clause[1][107] 	= partial_clause_prev[1][107] & 1'b1;
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & 1'b1;
			partial_clause[1][110] 	= partial_clause_prev[1][110] & 1'b1;
			partial_clause[1][111] 	= partial_clause_prev[1][111] & ~x[33];
			partial_clause[1][112] 	= partial_clause_prev[1][112] & 1'b1;
			partial_clause[1][113] 	= partial_clause_prev[1][113] & 1'b1;
			partial_clause[1][114] 	= partial_clause_prev[1][114] & 1'b1;
			partial_clause[1][115] 	= partial_clause_prev[1][115] & 1'b1;
			partial_clause[1][116] 	= partial_clause_prev[1][116] & x[2];
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & 1'b1;
			partial_clause[1][119] 	= partial_clause_prev[1][119] & 1'b1;
			partial_clause[1][120] 	= partial_clause_prev[1][120] & 1'b1;
			partial_clause[1][121] 	= partial_clause_prev[1][121] & 1'b1;
			partial_clause[1][122] 	= partial_clause_prev[1][122] & 1'b1;
			partial_clause[1][123] 	= partial_clause_prev[1][123] & 1'b1;
			partial_clause[1][124] 	= partial_clause_prev[1][124] & 1'b1;
			partial_clause[1][125] 	= partial_clause_prev[1][125] & 1'b1;
			partial_clause[1][126] 	= partial_clause_prev[1][126] & 1'b1;
			partial_clause[1][127] 	= partial_clause_prev[1][127] & ~x[34];
			partial_clause[1][128] 	= partial_clause_prev[1][128] & ~x[4];
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & ~x[2];
			partial_clause[1][131] 	= partial_clause_prev[1][131] & 1'b1;
			partial_clause[1][132] 	= partial_clause_prev[1][132] & 1'b1;
			partial_clause[1][133] 	= partial_clause_prev[1][133] & 1'b1;
			partial_clause[1][134] 	= partial_clause_prev[1][134] & 1'b1;
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & 1'b1;
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & 1'b1;
			partial_clause[1][139] 	= partial_clause_prev[1][139] & x[27];
			partial_clause[1][140] 	= partial_clause_prev[1][140] & 1'b1;
			partial_clause[1][141] 	= partial_clause_prev[1][141] & 1'b1;
			partial_clause[1][142] 	= partial_clause_prev[1][142] & x[4];
			partial_clause[1][143] 	= partial_clause_prev[1][143] & 1'b1;
			partial_clause[1][144] 	= partial_clause_prev[1][144] & 1'b1;
			partial_clause[1][145] 	= partial_clause_prev[1][145] & 1'b1;
			partial_clause[1][146] 	= partial_clause_prev[1][146] & 1'b1;
			partial_clause[1][147] 	= partial_clause_prev[1][147] & 1'b1;
			partial_clause[1][148] 	= partial_clause_prev[1][148] & 1'b1;
			partial_clause[1][149] 	= partial_clause_prev[1][149] & 1'b1;
			partial_clause[1][150] 	= partial_clause_prev[1][150] & 1'b1;
			partial_clause[1][151] 	= partial_clause_prev[1][151] & 1'b1;
			partial_clause[1][152] 	= partial_clause_prev[1][152] & 1'b1;
			partial_clause[1][153] 	= partial_clause_prev[1][153] & 1'b1;
			partial_clause[1][154] 	= partial_clause_prev[1][154] & 1'b1;
			partial_clause[1][155] 	= partial_clause_prev[1][155] & 1'b1;
			partial_clause[1][156] 	= partial_clause_prev[1][156] & 1'b1;
			partial_clause[1][157] 	= partial_clause_prev[1][157] & x[9];
			partial_clause[1][158] 	= partial_clause_prev[1][158] & x[1] & x[62];
			partial_clause[1][159] 	= partial_clause_prev[1][159] & 1'b1;
			partial_clause[1][160] 	= partial_clause_prev[1][160] & ~x[4] & ~x[44];
			partial_clause[1][161] 	= partial_clause_prev[1][161] & 1'b1;
			partial_clause[1][162] 	= partial_clause_prev[1][162] & 1'b1;
			partial_clause[1][163] 	= partial_clause_prev[1][163] & 1'b1;
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & 1'b1;
			partial_clause[1][166] 	= partial_clause_prev[1][166] & 1'b1;
			partial_clause[1][167] 	= partial_clause_prev[1][167] & x[11];
			partial_clause[1][168] 	= partial_clause_prev[1][168] & 1'b1;
			partial_clause[1][169] 	= partial_clause_prev[1][169] & 1'b1;
			partial_clause[1][170] 	= partial_clause_prev[1][170] & 1'b1;
			partial_clause[1][171] 	= partial_clause_prev[1][171] & 1'b1;
			partial_clause[1][172] 	= partial_clause_prev[1][172] & 1'b1;
			partial_clause[1][173] 	= partial_clause_prev[1][173] & 1'b1;
			partial_clause[1][174] 	= partial_clause_prev[1][174] & 1'b1;
			partial_clause[1][175] 	= partial_clause_prev[1][175] & 1'b1;
			partial_clause[1][176] 	= partial_clause_prev[1][176] & 1'b1;
			partial_clause[1][177] 	= partial_clause_prev[1][177] & 1'b1;
			partial_clause[1][178] 	= partial_clause_prev[1][178] & x[2];
			partial_clause[1][179] 	= partial_clause_prev[1][179] & 1'b1;
			partial_clause[1][180] 	= partial_clause_prev[1][180] & 1'b1;
			partial_clause[1][181] 	= partial_clause_prev[1][181] & 1'b1;
			partial_clause[1][182] 	= partial_clause_prev[1][182] & 1'b1;
			partial_clause[1][183] 	= partial_clause_prev[1][183] & 1'b1;
			partial_clause[1][184] 	= partial_clause_prev[1][184] & ~x[35];
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & 1'b1;
			partial_clause[1][187] 	= partial_clause_prev[1][187] & ~x[6] & x[9];
			partial_clause[1][188] 	= partial_clause_prev[1][188] & 1'b1;
			partial_clause[1][189] 	= partial_clause_prev[1][189] & 1'b1;
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & 1'b1;
			partial_clause[1][192] 	= partial_clause_prev[1][192] & 1'b1;
			partial_clause[1][193] 	= partial_clause_prev[1][193] & 1'b1;
			partial_clause[1][194] 	= partial_clause_prev[1][194] & 1'b1;
			partial_clause[1][195] 	= partial_clause_prev[1][195] & 1'b1;
			partial_clause[1][196] 	= partial_clause_prev[1][196] & 1'b1;
			partial_clause[1][197] 	= partial_clause_prev[1][197] & 1'b1;
			partial_clause[1][198] 	= partial_clause_prev[1][198] & 1'b1;
			partial_clause[1][199] 	= partial_clause_prev[1][199] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & x[4];
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & x[27];
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & x[16];
			partial_clause[2][7] 	= partial_clause_prev[2][7] & x[43];
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & x[31];
			partial_clause[2][11] 	= partial_clause_prev[2][11] & x[18];
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & x[55];
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & x[24];
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & x[12];
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & x[59];
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & ~x[10];
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & x[43];
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & x[16];
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & x[44];
			partial_clause[2][65] 	= partial_clause_prev[2][65] & x[8];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & x[41];
			partial_clause[2][69] 	= partial_clause_prev[2][69] & x[56];
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & x[16];
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & x[16];
			partial_clause[2][79] 	= partial_clause_prev[2][79] & x[0];
			partial_clause[2][80] 	= partial_clause_prev[2][80] & x[26];
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & x[44];
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & x[3];
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & x[25];
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & x[33];
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & x[5] & x[42];
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & x[13];
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			partial_clause[2][100] 	= partial_clause_prev[2][100] & ~x[42];
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & ~x[3];
			partial_clause[2][103] 	= partial_clause_prev[2][103] & 1'b1;
			partial_clause[2][104] 	= partial_clause_prev[2][104] & ~x[38];
			partial_clause[2][105] 	= partial_clause_prev[2][105] & ~x[40];
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & 1'b1;
			partial_clause[2][108] 	= partial_clause_prev[2][108] & 1'b1;
			partial_clause[2][109] 	= partial_clause_prev[2][109] & 1'b1;
			partial_clause[2][110] 	= partial_clause_prev[2][110] & 1'b1;
			partial_clause[2][111] 	= partial_clause_prev[2][111] & 1'b1;
			partial_clause[2][112] 	= partial_clause_prev[2][112] & 1'b1;
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & 1'b1;
			partial_clause[2][115] 	= partial_clause_prev[2][115] & 1'b1;
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & 1'b1;
			partial_clause[2][118] 	= partial_clause_prev[2][118] & ~x[12];
			partial_clause[2][119] 	= partial_clause_prev[2][119] & 1'b1;
			partial_clause[2][120] 	= partial_clause_prev[2][120] & 1'b1;
			partial_clause[2][121] 	= partial_clause_prev[2][121] & ~x[15] & ~x[59];
			partial_clause[2][122] 	= partial_clause_prev[2][122] & 1'b1;
			partial_clause[2][123] 	= partial_clause_prev[2][123] & 1'b1;
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & 1'b1;
			partial_clause[2][126] 	= partial_clause_prev[2][126] & 1'b1;
			partial_clause[2][127] 	= partial_clause_prev[2][127] & 1'b1;
			partial_clause[2][128] 	= partial_clause_prev[2][128] & 1'b1;
			partial_clause[2][129] 	= partial_clause_prev[2][129] & 1'b1;
			partial_clause[2][130] 	= partial_clause_prev[2][130] & 1'b1;
			partial_clause[2][131] 	= partial_clause_prev[2][131] & 1'b1;
			partial_clause[2][132] 	= partial_clause_prev[2][132] & 1'b1;
			partial_clause[2][133] 	= partial_clause_prev[2][133] & 1'b1;
			partial_clause[2][134] 	= partial_clause_prev[2][134] & 1'b1;
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & 1'b1;
			partial_clause[2][137] 	= partial_clause_prev[2][137] & 1'b1;
			partial_clause[2][138] 	= partial_clause_prev[2][138] & 1'b1;
			partial_clause[2][139] 	= partial_clause_prev[2][139] & 1'b1;
			partial_clause[2][140] 	= partial_clause_prev[2][140] & 1'b1;
			partial_clause[2][141] 	= partial_clause_prev[2][141] & 1'b1;
			partial_clause[2][142] 	= partial_clause_prev[2][142] & 1'b1;
			partial_clause[2][143] 	= partial_clause_prev[2][143] & 1'b1;
			partial_clause[2][144] 	= partial_clause_prev[2][144] & 1'b1;
			partial_clause[2][145] 	= partial_clause_prev[2][145] & ~x[2] & ~x[34];
			partial_clause[2][146] 	= partial_clause_prev[2][146] & 1'b1;
			partial_clause[2][147] 	= partial_clause_prev[2][147] & 1'b1;
			partial_clause[2][148] 	= partial_clause_prev[2][148] & ~x[4];
			partial_clause[2][149] 	= partial_clause_prev[2][149] & 1'b1;
			partial_clause[2][150] 	= partial_clause_prev[2][150] & ~x[34];
			partial_clause[2][151] 	= partial_clause_prev[2][151] & 1'b1;
			partial_clause[2][152] 	= partial_clause_prev[2][152] & 1'b1;
			partial_clause[2][153] 	= partial_clause_prev[2][153] & 1'b1;
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & ~x[41];
			partial_clause[2][156] 	= partial_clause_prev[2][156] & 1'b1;
			partial_clause[2][157] 	= partial_clause_prev[2][157] & 1'b1;
			partial_clause[2][158] 	= partial_clause_prev[2][158] & 1'b1;
			partial_clause[2][159] 	= partial_clause_prev[2][159] & 1'b1;
			partial_clause[2][160] 	= partial_clause_prev[2][160] & 1'b1;
			partial_clause[2][161] 	= partial_clause_prev[2][161] & ~x[11];
			partial_clause[2][162] 	= partial_clause_prev[2][162] & 1'b1;
			partial_clause[2][163] 	= partial_clause_prev[2][163] & 1'b1;
			partial_clause[2][164] 	= partial_clause_prev[2][164] & 1'b1;
			partial_clause[2][165] 	= partial_clause_prev[2][165] & 1'b1;
			partial_clause[2][166] 	= partial_clause_prev[2][166] & ~x[2] & ~x[4] & ~x[31] & ~x[60];
			partial_clause[2][167] 	= partial_clause_prev[2][167] & 1'b1;
			partial_clause[2][168] 	= partial_clause_prev[2][168] & ~x[0] & ~x[12];
			partial_clause[2][169] 	= partial_clause_prev[2][169] & 1'b1;
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & 1'b1;
			partial_clause[2][173] 	= partial_clause_prev[2][173] & 1'b1;
			partial_clause[2][174] 	= partial_clause_prev[2][174] & 1'b1;
			partial_clause[2][175] 	= partial_clause_prev[2][175] & 1'b1;
			partial_clause[2][176] 	= partial_clause_prev[2][176] & ~x[1] & ~x[43];
			partial_clause[2][177] 	= partial_clause_prev[2][177] & 1'b1;
			partial_clause[2][178] 	= partial_clause_prev[2][178] & ~x[42];
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & 1'b1;
			partial_clause[2][181] 	= partial_clause_prev[2][181] & ~x[15] & ~x[57];
			partial_clause[2][182] 	= partial_clause_prev[2][182] & 1'b1;
			partial_clause[2][183] 	= partial_clause_prev[2][183] & 1'b1;
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & 1'b1;
			partial_clause[2][186] 	= partial_clause_prev[2][186] & 1'b1;
			partial_clause[2][187] 	= partial_clause_prev[2][187] & 1'b1;
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & ~x[13];
			partial_clause[2][190] 	= partial_clause_prev[2][190] & ~x[5] & ~x[7];
			partial_clause[2][191] 	= partial_clause_prev[2][191] & 1'b1;
			partial_clause[2][192] 	= partial_clause_prev[2][192] & 1'b1;
			partial_clause[2][193] 	= partial_clause_prev[2][193] & ~x[32];
			partial_clause[2][194] 	= partial_clause_prev[2][194] & 1'b1;
			partial_clause[2][195] 	= partial_clause_prev[2][195] & ~x[3] & ~x[30];
			partial_clause[2][196] 	= partial_clause_prev[2][196] & ~x[2] & ~x[34];
			partial_clause[2][197] 	= partial_clause_prev[2][197] & 1'b1;
			partial_clause[2][198] 	= partial_clause_prev[2][198] & 1'b1;
			partial_clause[2][199] 	= partial_clause_prev[2][199] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & ~x[5];
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & ~x[7];
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & ~x[6];
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & x[52];
			partial_clause[3][24] 	= partial_clause_prev[3][24] & ~x[2];
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & ~x[4];
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & ~x[29] & ~x[30] & ~x[32] & ~x[33];
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & ~x[30];
			partial_clause[3][38] 	= partial_clause_prev[3][38] & ~x[5];
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & ~x[44];
			partial_clause[3][42] 	= partial_clause_prev[3][42] & x[9];
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & x[23];
			partial_clause[3][49] 	= partial_clause_prev[3][49] & ~x[31];
			partial_clause[3][50] 	= partial_clause_prev[3][50] & x[24];
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & ~x[1] & ~x[31] & ~x[33];
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & 1'b1;
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & ~x[1] & ~x[4];
			partial_clause[3][75] 	= partial_clause_prev[3][75] & x[24];
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & ~x[60] & ~x[62];
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & x[41];
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & x[51];
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & ~x[1] & ~x[32];
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			partial_clause[3][100] 	= partial_clause_prev[3][100] & 1'b1;
			partial_clause[3][101] 	= partial_clause_prev[3][101] & 1'b1;
			partial_clause[3][102] 	= partial_clause_prev[3][102] & ~x[9];
			partial_clause[3][103] 	= partial_clause_prev[3][103] & 1'b1;
			partial_clause[3][104] 	= partial_clause_prev[3][104] & 1'b1;
			partial_clause[3][105] 	= partial_clause_prev[3][105] & 1'b1;
			partial_clause[3][106] 	= partial_clause_prev[3][106] & 1'b1;
			partial_clause[3][107] 	= partial_clause_prev[3][107] & ~x[25] & x[32] & ~x[63];
			partial_clause[3][108] 	= partial_clause_prev[3][108] & x[29];
			partial_clause[3][109] 	= partial_clause_prev[3][109] & 1'b1;
			partial_clause[3][110] 	= partial_clause_prev[3][110] & x[62];
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & 1'b1;
			partial_clause[3][113] 	= partial_clause_prev[3][113] & ~x[27];
			partial_clause[3][114] 	= partial_clause_prev[3][114] & 1'b1;
			partial_clause[3][115] 	= partial_clause_prev[3][115] & 1'b1;
			partial_clause[3][116] 	= partial_clause_prev[3][116] & 1'b1;
			partial_clause[3][117] 	= partial_clause_prev[3][117] & 1'b1;
			partial_clause[3][118] 	= partial_clause_prev[3][118] & ~x[8];
			partial_clause[3][119] 	= partial_clause_prev[3][119] & 1'b1;
			partial_clause[3][120] 	= partial_clause_prev[3][120] & 1'b1;
			partial_clause[3][121] 	= partial_clause_prev[3][121] & 1'b1;
			partial_clause[3][122] 	= partial_clause_prev[3][122] & 1'b1;
			partial_clause[3][123] 	= partial_clause_prev[3][123] & x[3];
			partial_clause[3][124] 	= partial_clause_prev[3][124] & x[3];
			partial_clause[3][125] 	= partial_clause_prev[3][125] & 1'b1;
			partial_clause[3][126] 	= partial_clause_prev[3][126] & 1'b1;
			partial_clause[3][127] 	= partial_clause_prev[3][127] & 1'b1;
			partial_clause[3][128] 	= partial_clause_prev[3][128] & 1'b1;
			partial_clause[3][129] 	= partial_clause_prev[3][129] & 1'b1;
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & 1'b1;
			partial_clause[3][132] 	= partial_clause_prev[3][132] & x[44];
			partial_clause[3][133] 	= partial_clause_prev[3][133] & ~x[54];
			partial_clause[3][134] 	= partial_clause_prev[3][134] & 1'b1;
			partial_clause[3][135] 	= partial_clause_prev[3][135] & 1'b1;
			partial_clause[3][136] 	= partial_clause_prev[3][136] & 1'b1;
			partial_clause[3][137] 	= partial_clause_prev[3][137] & 1'b1;
			partial_clause[3][138] 	= partial_clause_prev[3][138] & x[5];
			partial_clause[3][139] 	= partial_clause_prev[3][139] & 1'b1;
			partial_clause[3][140] 	= partial_clause_prev[3][140] & 1'b1;
			partial_clause[3][141] 	= partial_clause_prev[3][141] & 1'b1;
			partial_clause[3][142] 	= partial_clause_prev[3][142] & x[58];
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & ~x[12] & x[34] & ~x[57];
			partial_clause[3][145] 	= partial_clause_prev[3][145] & ~x[9];
			partial_clause[3][146] 	= partial_clause_prev[3][146] & 1'b1;
			partial_clause[3][147] 	= partial_clause_prev[3][147] & 1'b1;
			partial_clause[3][148] 	= partial_clause_prev[3][148] & 1'b1;
			partial_clause[3][149] 	= partial_clause_prev[3][149] & ~x[14] & ~x[53];
			partial_clause[3][150] 	= partial_clause_prev[3][150] & 1'b1;
			partial_clause[3][151] 	= partial_clause_prev[3][151] & 1'b1;
			partial_clause[3][152] 	= partial_clause_prev[3][152] & x[60];
			partial_clause[3][153] 	= partial_clause_prev[3][153] & 1'b1;
			partial_clause[3][154] 	= partial_clause_prev[3][154] & 1'b1;
			partial_clause[3][155] 	= partial_clause_prev[3][155] & 1'b1;
			partial_clause[3][156] 	= partial_clause_prev[3][156] & ~x[37];
			partial_clause[3][157] 	= partial_clause_prev[3][157] & 1'b1;
			partial_clause[3][158] 	= partial_clause_prev[3][158] & 1'b1;
			partial_clause[3][159] 	= partial_clause_prev[3][159] & x[31];
			partial_clause[3][160] 	= partial_clause_prev[3][160] & x[5] & ~x[8];
			partial_clause[3][161] 	= partial_clause_prev[3][161] & 1'b1;
			partial_clause[3][162] 	= partial_clause_prev[3][162] & x[44];
			partial_clause[3][163] 	= partial_clause_prev[3][163] & 1'b1;
			partial_clause[3][164] 	= partial_clause_prev[3][164] & x[1];
			partial_clause[3][165] 	= partial_clause_prev[3][165] & 1'b1;
			partial_clause[3][166] 	= partial_clause_prev[3][166] & 1'b1;
			partial_clause[3][167] 	= partial_clause_prev[3][167] & x[60];
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & 1'b1;
			partial_clause[3][170] 	= partial_clause_prev[3][170] & 1'b1;
			partial_clause[3][171] 	= partial_clause_prev[3][171] & x[33];
			partial_clause[3][172] 	= partial_clause_prev[3][172] & 1'b1;
			partial_clause[3][173] 	= partial_clause_prev[3][173] & ~x[23];
			partial_clause[3][174] 	= partial_clause_prev[3][174] & x[0];
			partial_clause[3][175] 	= partial_clause_prev[3][175] & x[5] & x[32];
			partial_clause[3][176] 	= partial_clause_prev[3][176] & 1'b1;
			partial_clause[3][177] 	= partial_clause_prev[3][177] & ~x[14];
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & 1'b1;
			partial_clause[3][180] 	= partial_clause_prev[3][180] & 1'b1;
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & 1'b1;
			partial_clause[3][183] 	= partial_clause_prev[3][183] & 1'b1;
			partial_clause[3][184] 	= partial_clause_prev[3][184] & 1'b1;
			partial_clause[3][185] 	= partial_clause_prev[3][185] & 1'b1;
			partial_clause[3][186] 	= partial_clause_prev[3][186] & ~x[42];
			partial_clause[3][187] 	= partial_clause_prev[3][187] & 1'b1;
			partial_clause[3][188] 	= partial_clause_prev[3][188] & 1'b1;
			partial_clause[3][189] 	= partial_clause_prev[3][189] & x[4] & x[59];
			partial_clause[3][190] 	= partial_clause_prev[3][190] & 1'b1;
			partial_clause[3][191] 	= partial_clause_prev[3][191] & 1'b1;
			partial_clause[3][192] 	= partial_clause_prev[3][192] & 1'b1;
			partial_clause[3][193] 	= partial_clause_prev[3][193] & 1'b1;
			partial_clause[3][194] 	= partial_clause_prev[3][194] & ~x[41];
			partial_clause[3][195] 	= partial_clause_prev[3][195] & 1'b1;
			partial_clause[3][196] 	= partial_clause_prev[3][196] & 1'b1;
			partial_clause[3][197] 	= partial_clause_prev[3][197] & x[16];
			partial_clause[3][198] 	= partial_clause_prev[3][198] & x[30];
			partial_clause[3][199] 	= partial_clause_prev[3][199] & ~x[51];
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & ~x[31];
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & ~x[12];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & ~x[60];
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & ~x[30] & ~x[56];
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & ~x[11];
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & ~x[61];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[40];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & ~x[38];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & ~x[32];
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[31];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & ~x[30] & ~x[32];
			partial_clause[4][51] 	= partial_clause_prev[4][51] & x[49];
			partial_clause[4][52] 	= partial_clause_prev[4][52] & ~x[32];
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & ~x[32];
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & ~x[62];
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & ~x[61];
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & ~x[27];
			partial_clause[4][80] 	= partial_clause_prev[4][80] & ~x[41];
			partial_clause[4][81] 	= partial_clause_prev[4][81] & ~x[40];
			partial_clause[4][82] 	= partial_clause_prev[4][82] & ~x[58];
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & ~x[61];
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & ~x[55];
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & ~x[28];
			partial_clause[4][100] 	= partial_clause_prev[4][100] & 1'b1;
			partial_clause[4][101] 	= partial_clause_prev[4][101] & 1'b1;
			partial_clause[4][102] 	= partial_clause_prev[4][102] & ~x[5];
			partial_clause[4][103] 	= partial_clause_prev[4][103] & 1'b1;
			partial_clause[4][104] 	= partial_clause_prev[4][104] & 1'b1;
			partial_clause[4][105] 	= partial_clause_prev[4][105] & 1'b1;
			partial_clause[4][106] 	= partial_clause_prev[4][106] & 1'b1;
			partial_clause[4][107] 	= partial_clause_prev[4][107] & ~x[5];
			partial_clause[4][108] 	= partial_clause_prev[4][108] & 1'b1;
			partial_clause[4][109] 	= partial_clause_prev[4][109] & 1'b1;
			partial_clause[4][110] 	= partial_clause_prev[4][110] & 1'b1;
			partial_clause[4][111] 	= partial_clause_prev[4][111] & 1'b1;
			partial_clause[4][112] 	= partial_clause_prev[4][112] & 1'b1;
			partial_clause[4][113] 	= partial_clause_prev[4][113] & x[60] & x[61];
			partial_clause[4][114] 	= partial_clause_prev[4][114] & 1'b1;
			partial_clause[4][115] 	= partial_clause_prev[4][115] & 1'b1;
			partial_clause[4][116] 	= partial_clause_prev[4][116] & x[30];
			partial_clause[4][117] 	= partial_clause_prev[4][117] & 1'b1;
			partial_clause[4][118] 	= partial_clause_prev[4][118] & x[56];
			partial_clause[4][119] 	= partial_clause_prev[4][119] & x[60];
			partial_clause[4][120] 	= partial_clause_prev[4][120] & 1'b1;
			partial_clause[4][121] 	= partial_clause_prev[4][121] & ~x[45];
			partial_clause[4][122] 	= partial_clause_prev[4][122] & 1'b1;
			partial_clause[4][123] 	= partial_clause_prev[4][123] & 1'b1;
			partial_clause[4][124] 	= partial_clause_prev[4][124] & 1'b1;
			partial_clause[4][125] 	= partial_clause_prev[4][125] & 1'b1;
			partial_clause[4][126] 	= partial_clause_prev[4][126] & 1'b1;
			partial_clause[4][127] 	= partial_clause_prev[4][127] & 1'b1;
			partial_clause[4][128] 	= partial_clause_prev[4][128] & x[30] & x[60];
			partial_clause[4][129] 	= partial_clause_prev[4][129] & 1'b1;
			partial_clause[4][130] 	= partial_clause_prev[4][130] & 1'b1;
			partial_clause[4][131] 	= partial_clause_prev[4][131] & 1'b1;
			partial_clause[4][132] 	= partial_clause_prev[4][132] & 1'b1;
			partial_clause[4][133] 	= partial_clause_prev[4][133] & 1'b1;
			partial_clause[4][134] 	= partial_clause_prev[4][134] & 1'b1;
			partial_clause[4][135] 	= partial_clause_prev[4][135] & 1'b1;
			partial_clause[4][136] 	= partial_clause_prev[4][136] & 1'b1;
			partial_clause[4][137] 	= partial_clause_prev[4][137] & 1'b1;
			partial_clause[4][138] 	= partial_clause_prev[4][138] & 1'b1;
			partial_clause[4][139] 	= partial_clause_prev[4][139] & 1'b1;
			partial_clause[4][140] 	= partial_clause_prev[4][140] & 1'b1;
			partial_clause[4][141] 	= partial_clause_prev[4][141] & x[42];
			partial_clause[4][142] 	= partial_clause_prev[4][142] & 1'b1;
			partial_clause[4][143] 	= partial_clause_prev[4][143] & 1'b1;
			partial_clause[4][144] 	= partial_clause_prev[4][144] & 1'b1;
			partial_clause[4][145] 	= partial_clause_prev[4][145] & 1'b1;
			partial_clause[4][146] 	= partial_clause_prev[4][146] & 1'b1;
			partial_clause[4][147] 	= partial_clause_prev[4][147] & 1'b1;
			partial_clause[4][148] 	= partial_clause_prev[4][148] & 1'b1;
			partial_clause[4][149] 	= partial_clause_prev[4][149] & 1'b1;
			partial_clause[4][150] 	= partial_clause_prev[4][150] & 1'b1;
			partial_clause[4][151] 	= partial_clause_prev[4][151] & 1'b1;
			partial_clause[4][152] 	= partial_clause_prev[4][152] & x[56];
			partial_clause[4][153] 	= partial_clause_prev[4][153] & 1'b1;
			partial_clause[4][154] 	= partial_clause_prev[4][154] & 1'b1;
			partial_clause[4][155] 	= partial_clause_prev[4][155] & 1'b1;
			partial_clause[4][156] 	= partial_clause_prev[4][156] & 1'b1;
			partial_clause[4][157] 	= partial_clause_prev[4][157] & 1'b1;
			partial_clause[4][158] 	= partial_clause_prev[4][158] & 1'b1;
			partial_clause[4][159] 	= partial_clause_prev[4][159] & 1'b1;
			partial_clause[4][160] 	= partial_clause_prev[4][160] & 1'b1;
			partial_clause[4][161] 	= partial_clause_prev[4][161] & 1'b1;
			partial_clause[4][162] 	= partial_clause_prev[4][162] & 1'b1;
			partial_clause[4][163] 	= partial_clause_prev[4][163] & x[59];
			partial_clause[4][164] 	= partial_clause_prev[4][164] & 1'b1;
			partial_clause[4][165] 	= partial_clause_prev[4][165] & 1'b1;
			partial_clause[4][166] 	= partial_clause_prev[4][166] & 1'b1;
			partial_clause[4][167] 	= partial_clause_prev[4][167] & 1'b1;
			partial_clause[4][168] 	= partial_clause_prev[4][168] & 1'b1;
			partial_clause[4][169] 	= partial_clause_prev[4][169] & 1'b1;
			partial_clause[4][170] 	= partial_clause_prev[4][170] & 1'b1;
			partial_clause[4][171] 	= partial_clause_prev[4][171] & 1'b1;
			partial_clause[4][172] 	= partial_clause_prev[4][172] & 1'b1;
			partial_clause[4][173] 	= partial_clause_prev[4][173] & 1'b1;
			partial_clause[4][174] 	= partial_clause_prev[4][174] & 1'b1;
			partial_clause[4][175] 	= partial_clause_prev[4][175] & 1'b1;
			partial_clause[4][176] 	= partial_clause_prev[4][176] & 1'b1;
			partial_clause[4][177] 	= partial_clause_prev[4][177] & 1'b1;
			partial_clause[4][178] 	= partial_clause_prev[4][178] & 1'b1;
			partial_clause[4][179] 	= partial_clause_prev[4][179] & 1'b1;
			partial_clause[4][180] 	= partial_clause_prev[4][180] & 1'b1;
			partial_clause[4][181] 	= partial_clause_prev[4][181] & 1'b1;
			partial_clause[4][182] 	= partial_clause_prev[4][182] & 1'b1;
			partial_clause[4][183] 	= partial_clause_prev[4][183] & 1'b1;
			partial_clause[4][184] 	= partial_clause_prev[4][184] & 1'b1;
			partial_clause[4][185] 	= partial_clause_prev[4][185] & x[29] & x[58];
			partial_clause[4][186] 	= partial_clause_prev[4][186] & 1'b1;
			partial_clause[4][187] 	= partial_clause_prev[4][187] & 1'b1;
			partial_clause[4][188] 	= partial_clause_prev[4][188] & x[58];
			partial_clause[4][189] 	= partial_clause_prev[4][189] & 1'b1;
			partial_clause[4][190] 	= partial_clause_prev[4][190] & 1'b1;
			partial_clause[4][191] 	= partial_clause_prev[4][191] & 1'b1;
			partial_clause[4][192] 	= partial_clause_prev[4][192] & x[39];
			partial_clause[4][193] 	= partial_clause_prev[4][193] & 1'b1;
			partial_clause[4][194] 	= partial_clause_prev[4][194] & x[60] & x[63];
			partial_clause[4][195] 	= partial_clause_prev[4][195] & 1'b1;
			partial_clause[4][196] 	= partial_clause_prev[4][196] & 1'b1;
			partial_clause[4][197] 	= partial_clause_prev[4][197] & 1'b1;
			partial_clause[4][198] 	= partial_clause_prev[4][198] & x[31];
			partial_clause[4][199] 	= partial_clause_prev[4][199] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & ~x[5];
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & ~x[8];
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & ~x[35];
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & ~x[2] & ~x[3];
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & ~x[33];
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & ~x[4];
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & ~x[4];
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & x[27];
			partial_clause[5][69] 	= partial_clause_prev[5][69] & ~x[0] & ~x[3] & ~x[5];
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & x[56];
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			partial_clause[5][100] 	= partial_clause_prev[5][100] & 1'b1;
			partial_clause[5][101] 	= partial_clause_prev[5][101] & 1'b1;
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & 1'b1;
			partial_clause[5][104] 	= partial_clause_prev[5][104] & 1'b1;
			partial_clause[5][105] 	= partial_clause_prev[5][105] & 1'b1;
			partial_clause[5][106] 	= partial_clause_prev[5][106] & 1'b1;
			partial_clause[5][107] 	= partial_clause_prev[5][107] & x[2];
			partial_clause[5][108] 	= partial_clause_prev[5][108] & 1'b1;
			partial_clause[5][109] 	= partial_clause_prev[5][109] & 1'b1;
			partial_clause[5][110] 	= partial_clause_prev[5][110] & 1'b1;
			partial_clause[5][111] 	= partial_clause_prev[5][111] & 1'b1;
			partial_clause[5][112] 	= partial_clause_prev[5][112] & 1'b1;
			partial_clause[5][113] 	= partial_clause_prev[5][113] & 1'b1;
			partial_clause[5][114] 	= partial_clause_prev[5][114] & 1'b1;
			partial_clause[5][115] 	= partial_clause_prev[5][115] & 1'b1;
			partial_clause[5][116] 	= partial_clause_prev[5][116] & 1'b1;
			partial_clause[5][117] 	= partial_clause_prev[5][117] & 1'b1;
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & 1'b1;
			partial_clause[5][120] 	= partial_clause_prev[5][120] & 1'b1;
			partial_clause[5][121] 	= partial_clause_prev[5][121] & 1'b1;
			partial_clause[5][122] 	= partial_clause_prev[5][122] & 1'b1;
			partial_clause[5][123] 	= partial_clause_prev[5][123] & 1'b1;
			partial_clause[5][124] 	= partial_clause_prev[5][124] & 1'b1;
			partial_clause[5][125] 	= partial_clause_prev[5][125] & 1'b1;
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & ~x[24] & ~x[26] & ~x[53];
			partial_clause[5][128] 	= partial_clause_prev[5][128] & x[3];
			partial_clause[5][129] 	= partial_clause_prev[5][129] & 1'b1;
			partial_clause[5][130] 	= partial_clause_prev[5][130] & 1'b1;
			partial_clause[5][131] 	= partial_clause_prev[5][131] & 1'b1;
			partial_clause[5][132] 	= partial_clause_prev[5][132] & ~x[57];
			partial_clause[5][133] 	= partial_clause_prev[5][133] & 1'b1;
			partial_clause[5][134] 	= partial_clause_prev[5][134] & x[29];
			partial_clause[5][135] 	= partial_clause_prev[5][135] & 1'b1;
			partial_clause[5][136] 	= partial_clause_prev[5][136] & 1'b1;
			partial_clause[5][137] 	= partial_clause_prev[5][137] & 1'b1;
			partial_clause[5][138] 	= partial_clause_prev[5][138] & 1'b1;
			partial_clause[5][139] 	= partial_clause_prev[5][139] & 1'b1;
			partial_clause[5][140] 	= partial_clause_prev[5][140] & 1'b1;
			partial_clause[5][141] 	= partial_clause_prev[5][141] & 1'b1;
			partial_clause[5][142] 	= partial_clause_prev[5][142] & 1'b1;
			partial_clause[5][143] 	= partial_clause_prev[5][143] & 1'b1;
			partial_clause[5][144] 	= partial_clause_prev[5][144] & 1'b1;
			partial_clause[5][145] 	= partial_clause_prev[5][145] & 1'b1;
			partial_clause[5][146] 	= partial_clause_prev[5][146] & x[29];
			partial_clause[5][147] 	= partial_clause_prev[5][147] & 1'b1;
			partial_clause[5][148] 	= partial_clause_prev[5][148] & 1'b1;
			partial_clause[5][149] 	= partial_clause_prev[5][149] & 1'b1;
			partial_clause[5][150] 	= partial_clause_prev[5][150] & 1'b1;
			partial_clause[5][151] 	= partial_clause_prev[5][151] & 1'b1;
			partial_clause[5][152] 	= partial_clause_prev[5][152] & 1'b1;
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & 1'b1;
			partial_clause[5][155] 	= partial_clause_prev[5][155] & 1'b1;
			partial_clause[5][156] 	= partial_clause_prev[5][156] & 1'b1;
			partial_clause[5][157] 	= partial_clause_prev[5][157] & 1'b1;
			partial_clause[5][158] 	= partial_clause_prev[5][158] & 1'b1;
			partial_clause[5][159] 	= partial_clause_prev[5][159] & 1'b1;
			partial_clause[5][160] 	= partial_clause_prev[5][160] & 1'b1;
			partial_clause[5][161] 	= partial_clause_prev[5][161] & 1'b1;
			partial_clause[5][162] 	= partial_clause_prev[5][162] & x[0];
			partial_clause[5][163] 	= partial_clause_prev[5][163] & 1'b1;
			partial_clause[5][164] 	= partial_clause_prev[5][164] & 1'b1;
			partial_clause[5][165] 	= partial_clause_prev[5][165] & x[2] & x[30];
			partial_clause[5][166] 	= partial_clause_prev[5][166] & 1'b1;
			partial_clause[5][167] 	= partial_clause_prev[5][167] & 1'b1;
			partial_clause[5][168] 	= partial_clause_prev[5][168] & 1'b1;
			partial_clause[5][169] 	= partial_clause_prev[5][169] & 1'b1;
			partial_clause[5][170] 	= partial_clause_prev[5][170] & 1'b1;
			partial_clause[5][171] 	= partial_clause_prev[5][171] & 1'b1;
			partial_clause[5][172] 	= partial_clause_prev[5][172] & 1'b1;
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & 1'b1;
			partial_clause[5][175] 	= partial_clause_prev[5][175] & 1'b1;
			partial_clause[5][176] 	= partial_clause_prev[5][176] & 1'b1;
			partial_clause[5][177] 	= partial_clause_prev[5][177] & 1'b1;
			partial_clause[5][178] 	= partial_clause_prev[5][178] & 1'b1;
			partial_clause[5][179] 	= partial_clause_prev[5][179] & 1'b1;
			partial_clause[5][180] 	= partial_clause_prev[5][180] & 1'b1;
			partial_clause[5][181] 	= partial_clause_prev[5][181] & 1'b1;
			partial_clause[5][182] 	= partial_clause_prev[5][182] & 1'b1;
			partial_clause[5][183] 	= partial_clause_prev[5][183] & 1'b1;
			partial_clause[5][184] 	= partial_clause_prev[5][184] & 1'b1;
			partial_clause[5][185] 	= partial_clause_prev[5][185] & 1'b1;
			partial_clause[5][186] 	= partial_clause_prev[5][186] & 1'b1;
			partial_clause[5][187] 	= partial_clause_prev[5][187] & 1'b1;
			partial_clause[5][188] 	= partial_clause_prev[5][188] & 1'b1;
			partial_clause[5][189] 	= partial_clause_prev[5][189] & ~x[58];
			partial_clause[5][190] 	= partial_clause_prev[5][190] & 1'b1;
			partial_clause[5][191] 	= partial_clause_prev[5][191] & 1'b1;
			partial_clause[5][192] 	= partial_clause_prev[5][192] & 1'b1;
			partial_clause[5][193] 	= partial_clause_prev[5][193] & x[5];
			partial_clause[5][194] 	= partial_clause_prev[5][194] & 1'b1;
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & 1'b1;
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & 1'b1;
			partial_clause[5][199] 	= partial_clause_prev[5][199] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & ~x[14];
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & x[62];
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & x[3];
			partial_clause[6][21] 	= partial_clause_prev[6][21] & x[30];
			partial_clause[6][22] 	= partial_clause_prev[6][22] & x[59];
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & x[5];
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & x[62];
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & x[30];
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & x[3];
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & x[58];
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & x[62];
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & x[63];
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & x[3];
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & x[63];
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			partial_clause[6][100] 	= partial_clause_prev[6][100] & ~x[36];
			partial_clause[6][101] 	= partial_clause_prev[6][101] & 1'b1;
			partial_clause[6][102] 	= partial_clause_prev[6][102] & 1'b1;
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & 1'b1;
			partial_clause[6][105] 	= partial_clause_prev[6][105] & x[43];
			partial_clause[6][106] 	= partial_clause_prev[6][106] & 1'b1;
			partial_clause[6][107] 	= partial_clause_prev[6][107] & 1'b1;
			partial_clause[6][108] 	= partial_clause_prev[6][108] & 1'b1;
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & 1'b1;
			partial_clause[6][111] 	= partial_clause_prev[6][111] & ~x[0] & ~x[2] & ~x[20];
			partial_clause[6][112] 	= partial_clause_prev[6][112] & ~x[1];
			partial_clause[6][113] 	= partial_clause_prev[6][113] & 1'b1;
			partial_clause[6][114] 	= partial_clause_prev[6][114] & 1'b1;
			partial_clause[6][115] 	= partial_clause_prev[6][115] & 1'b1;
			partial_clause[6][116] 	= partial_clause_prev[6][116] & 1'b1;
			partial_clause[6][117] 	= partial_clause_prev[6][117] & ~x[60];
			partial_clause[6][118] 	= partial_clause_prev[6][118] & 1'b1;
			partial_clause[6][119] 	= partial_clause_prev[6][119] & 1'b1;
			partial_clause[6][120] 	= partial_clause_prev[6][120] & 1'b1;
			partial_clause[6][121] 	= partial_clause_prev[6][121] & x[56];
			partial_clause[6][122] 	= partial_clause_prev[6][122] & 1'b1;
			partial_clause[6][123] 	= partial_clause_prev[6][123] & ~x[36];
			partial_clause[6][124] 	= partial_clause_prev[6][124] & 1'b1;
			partial_clause[6][125] 	= partial_clause_prev[6][125] & 1'b1;
			partial_clause[6][126] 	= partial_clause_prev[6][126] & 1'b1;
			partial_clause[6][127] 	= partial_clause_prev[6][127] & 1'b1;
			partial_clause[6][128] 	= partial_clause_prev[6][128] & 1'b1;
			partial_clause[6][129] 	= partial_clause_prev[6][129] & 1'b1;
			partial_clause[6][130] 	= partial_clause_prev[6][130] & 1'b1;
			partial_clause[6][131] 	= partial_clause_prev[6][131] & 1'b1;
			partial_clause[6][132] 	= partial_clause_prev[6][132] & 1'b1;
			partial_clause[6][133] 	= partial_clause_prev[6][133] & 1'b1;
			partial_clause[6][134] 	= partial_clause_prev[6][134] & 1'b1;
			partial_clause[6][135] 	= partial_clause_prev[6][135] & ~x[29];
			partial_clause[6][136] 	= partial_clause_prev[6][136] & 1'b1;
			partial_clause[6][137] 	= partial_clause_prev[6][137] & 1'b1;
			partial_clause[6][138] 	= partial_clause_prev[6][138] & 1'b1;
			partial_clause[6][139] 	= partial_clause_prev[6][139] & 1'b1;
			partial_clause[6][140] 	= partial_clause_prev[6][140] & 1'b1;
			partial_clause[6][141] 	= partial_clause_prev[6][141] & ~x[31] & ~x[56];
			partial_clause[6][142] 	= partial_clause_prev[6][142] & 1'b1;
			partial_clause[6][143] 	= partial_clause_prev[6][143] & 1'b1;
			partial_clause[6][144] 	= partial_clause_prev[6][144] & 1'b1;
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & 1'b1;
			partial_clause[6][147] 	= partial_clause_prev[6][147] & 1'b1;
			partial_clause[6][148] 	= partial_clause_prev[6][148] & 1'b1;
			partial_clause[6][149] 	= partial_clause_prev[6][149] & x[52];
			partial_clause[6][150] 	= partial_clause_prev[6][150] & ~x[3] & ~x[4] & ~x[28] & ~x[30];
			partial_clause[6][151] 	= partial_clause_prev[6][151] & 1'b1;
			partial_clause[6][152] 	= partial_clause_prev[6][152] & ~x[33];
			partial_clause[6][153] 	= partial_clause_prev[6][153] & 1'b1;
			partial_clause[6][154] 	= partial_clause_prev[6][154] & 1'b1;
			partial_clause[6][155] 	= partial_clause_prev[6][155] & x[26];
			partial_clause[6][156] 	= partial_clause_prev[6][156] & 1'b1;
			partial_clause[6][157] 	= partial_clause_prev[6][157] & ~x[1] & ~x[3];
			partial_clause[6][158] 	= partial_clause_prev[6][158] & 1'b1;
			partial_clause[6][159] 	= partial_clause_prev[6][159] & 1'b1;
			partial_clause[6][160] 	= partial_clause_prev[6][160] & 1'b1;
			partial_clause[6][161] 	= partial_clause_prev[6][161] & 1'b1;
			partial_clause[6][162] 	= partial_clause_prev[6][162] & 1'b1;
			partial_clause[6][163] 	= partial_clause_prev[6][163] & ~x[33] & ~x[60];
			partial_clause[6][164] 	= partial_clause_prev[6][164] & 1'b1;
			partial_clause[6][165] 	= partial_clause_prev[6][165] & 1'b1;
			partial_clause[6][166] 	= partial_clause_prev[6][166] & 1'b1;
			partial_clause[6][167] 	= partial_clause_prev[6][167] & 1'b1;
			partial_clause[6][168] 	= partial_clause_prev[6][168] & 1'b1;
			partial_clause[6][169] 	= partial_clause_prev[6][169] & 1'b1;
			partial_clause[6][170] 	= partial_clause_prev[6][170] & 1'b1;
			partial_clause[6][171] 	= partial_clause_prev[6][171] & ~x[32] & ~x[59];
			partial_clause[6][172] 	= partial_clause_prev[6][172] & 1'b1;
			partial_clause[6][173] 	= partial_clause_prev[6][173] & 1'b1;
			partial_clause[6][174] 	= partial_clause_prev[6][174] & ~x[29];
			partial_clause[6][175] 	= partial_clause_prev[6][175] & 1'b1;
			partial_clause[6][176] 	= partial_clause_prev[6][176] & 1'b1;
			partial_clause[6][177] 	= partial_clause_prev[6][177] & ~x[32] & ~x[59];
			partial_clause[6][178] 	= partial_clause_prev[6][178] & 1'b1;
			partial_clause[6][179] 	= partial_clause_prev[6][179] & 1'b1;
			partial_clause[6][180] 	= partial_clause_prev[6][180] & 1'b1;
			partial_clause[6][181] 	= partial_clause_prev[6][181] & ~x[62];
			partial_clause[6][182] 	= partial_clause_prev[6][182] & ~x[29];
			partial_clause[6][183] 	= partial_clause_prev[6][183] & 1'b1;
			partial_clause[6][184] 	= partial_clause_prev[6][184] & 1'b1;
			partial_clause[6][185] 	= partial_clause_prev[6][185] & 1'b1;
			partial_clause[6][186] 	= partial_clause_prev[6][186] & 1'b1;
			partial_clause[6][187] 	= partial_clause_prev[6][187] & 1'b1;
			partial_clause[6][188] 	= partial_clause_prev[6][188] & 1'b1;
			partial_clause[6][189] 	= partial_clause_prev[6][189] & ~x[4] & ~x[28] & ~x[30];
			partial_clause[6][190] 	= partial_clause_prev[6][190] & ~x[32] & ~x[57] & ~x[59];
			partial_clause[6][191] 	= partial_clause_prev[6][191] & 1'b1;
			partial_clause[6][192] 	= partial_clause_prev[6][192] & 1'b1;
			partial_clause[6][193] 	= partial_clause_prev[6][193] & 1'b1;
			partial_clause[6][194] 	= partial_clause_prev[6][194] & 1'b1;
			partial_clause[6][195] 	= partial_clause_prev[6][195] & 1'b1;
			partial_clause[6][196] 	= partial_clause_prev[6][196] & 1'b1;
			partial_clause[6][197] 	= partial_clause_prev[6][197] & 1'b1;
			partial_clause[6][198] 	= partial_clause_prev[6][198] & 1'b1;
			partial_clause[6][199] 	= partial_clause_prev[6][199] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & ~x[57];
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & ~x[2];
			partial_clause[7][9] 	= partial_clause_prev[7][9] & ~x[31];
			partial_clause[7][10] 	= partial_clause_prev[7][10] & x[32];
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & ~x[30];
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & ~x[39];
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & ~x[30];
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & ~x[10];
			partial_clause[7][40] 	= partial_clause_prev[7][40] & ~x[13];
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & ~x[14];
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & x[20];
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & ~x[2];
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & ~x[2] & ~x[58];
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & ~x[39] & ~x[40];
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & ~x[53];
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & ~x[39];
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & ~x[1];
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			partial_clause[7][100] 	= partial_clause_prev[7][100] & 1'b1;
			partial_clause[7][101] 	= partial_clause_prev[7][101] & 1'b1;
			partial_clause[7][102] 	= partial_clause_prev[7][102] & 1'b1;
			partial_clause[7][103] 	= partial_clause_prev[7][103] & 1'b1;
			partial_clause[7][104] 	= partial_clause_prev[7][104] & 1'b1;
			partial_clause[7][105] 	= partial_clause_prev[7][105] & 1'b1;
			partial_clause[7][106] 	= partial_clause_prev[7][106] & 1'b1;
			partial_clause[7][107] 	= partial_clause_prev[7][107] & 1'b1;
			partial_clause[7][108] 	= partial_clause_prev[7][108] & 1'b1;
			partial_clause[7][109] 	= partial_clause_prev[7][109] & ~x[50];
			partial_clause[7][110] 	= partial_clause_prev[7][110] & 1'b1;
			partial_clause[7][111] 	= partial_clause_prev[7][111] & 1'b1;
			partial_clause[7][112] 	= partial_clause_prev[7][112] & x[26];
			partial_clause[7][113] 	= partial_clause_prev[7][113] & 1'b1;
			partial_clause[7][114] 	= partial_clause_prev[7][114] & 1'b1;
			partial_clause[7][115] 	= partial_clause_prev[7][115] & 1'b1;
			partial_clause[7][116] 	= partial_clause_prev[7][116] & 1'b1;
			partial_clause[7][117] 	= partial_clause_prev[7][117] & x[41];
			partial_clause[7][118] 	= partial_clause_prev[7][118] & 1'b1;
			partial_clause[7][119] 	= partial_clause_prev[7][119] & x[2];
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & 1'b1;
			partial_clause[7][123] 	= partial_clause_prev[7][123] & x[25];
			partial_clause[7][124] 	= partial_clause_prev[7][124] & 1'b1;
			partial_clause[7][125] 	= partial_clause_prev[7][125] & 1'b1;
			partial_clause[7][126] 	= partial_clause_prev[7][126] & 1'b1;
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & 1'b1;
			partial_clause[7][129] 	= partial_clause_prev[7][129] & x[8];
			partial_clause[7][130] 	= partial_clause_prev[7][130] & 1'b1;
			partial_clause[7][131] 	= partial_clause_prev[7][131] & 1'b1;
			partial_clause[7][132] 	= partial_clause_prev[7][132] & 1'b1;
			partial_clause[7][133] 	= partial_clause_prev[7][133] & 1'b1;
			partial_clause[7][134] 	= partial_clause_prev[7][134] & x[41];
			partial_clause[7][135] 	= partial_clause_prev[7][135] & 1'b1;
			partial_clause[7][136] 	= partial_clause_prev[7][136] & 1'b1;
			partial_clause[7][137] 	= partial_clause_prev[7][137] & 1'b1;
			partial_clause[7][138] 	= partial_clause_prev[7][138] & x[2];
			partial_clause[7][139] 	= partial_clause_prev[7][139] & 1'b1;
			partial_clause[7][140] 	= partial_clause_prev[7][140] & 1'b1;
			partial_clause[7][141] 	= partial_clause_prev[7][141] & 1'b1;
			partial_clause[7][142] 	= partial_clause_prev[7][142] & 1'b1;
			partial_clause[7][143] 	= partial_clause_prev[7][143] & x[27];
			partial_clause[7][144] 	= partial_clause_prev[7][144] & 1'b1;
			partial_clause[7][145] 	= partial_clause_prev[7][145] & 1'b1;
			partial_clause[7][146] 	= partial_clause_prev[7][146] & 1'b1;
			partial_clause[7][147] 	= partial_clause_prev[7][147] & 1'b1;
			partial_clause[7][148] 	= partial_clause_prev[7][148] & 1'b1;
			partial_clause[7][149] 	= partial_clause_prev[7][149] & 1'b1;
			partial_clause[7][150] 	= partial_clause_prev[7][150] & 1'b1;
			partial_clause[7][151] 	= partial_clause_prev[7][151] & 1'b1;
			partial_clause[7][152] 	= partial_clause_prev[7][152] & 1'b1;
			partial_clause[7][153] 	= partial_clause_prev[7][153] & 1'b1;
			partial_clause[7][154] 	= partial_clause_prev[7][154] & 1'b1;
			partial_clause[7][155] 	= partial_clause_prev[7][155] & 1'b1;
			partial_clause[7][156] 	= partial_clause_prev[7][156] & 1'b1;
			partial_clause[7][157] 	= partial_clause_prev[7][157] & 1'b1;
			partial_clause[7][158] 	= partial_clause_prev[7][158] & 1'b1;
			partial_clause[7][159] 	= partial_clause_prev[7][159] & 1'b1;
			partial_clause[7][160] 	= partial_clause_prev[7][160] & 1'b1;
			partial_clause[7][161] 	= partial_clause_prev[7][161] & 1'b1;
			partial_clause[7][162] 	= partial_clause_prev[7][162] & 1'b1;
			partial_clause[7][163] 	= partial_clause_prev[7][163] & 1'b1;
			partial_clause[7][164] 	= partial_clause_prev[7][164] & 1'b1;
			partial_clause[7][165] 	= partial_clause_prev[7][165] & 1'b1;
			partial_clause[7][166] 	= partial_clause_prev[7][166] & 1'b1;
			partial_clause[7][167] 	= partial_clause_prev[7][167] & 1'b1;
			partial_clause[7][168] 	= partial_clause_prev[7][168] & 1'b1;
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & 1'b1;
			partial_clause[7][171] 	= partial_clause_prev[7][171] & 1'b1;
			partial_clause[7][172] 	= partial_clause_prev[7][172] & 1'b1;
			partial_clause[7][173] 	= partial_clause_prev[7][173] & 1'b1;
			partial_clause[7][174] 	= partial_clause_prev[7][174] & 1'b1;
			partial_clause[7][175] 	= partial_clause_prev[7][175] & x[57];
			partial_clause[7][176] 	= partial_clause_prev[7][176] & 1'b1;
			partial_clause[7][177] 	= partial_clause_prev[7][177] & x[27];
			partial_clause[7][178] 	= partial_clause_prev[7][178] & 1'b1;
			partial_clause[7][179] 	= partial_clause_prev[7][179] & 1'b1;
			partial_clause[7][180] 	= partial_clause_prev[7][180] & 1'b1;
			partial_clause[7][181] 	= partial_clause_prev[7][181] & 1'b1;
			partial_clause[7][182] 	= partial_clause_prev[7][182] & x[0];
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & x[25];
			partial_clause[7][185] 	= partial_clause_prev[7][185] & 1'b1;
			partial_clause[7][186] 	= partial_clause_prev[7][186] & 1'b1;
			partial_clause[7][187] 	= partial_clause_prev[7][187] & x[36];
			partial_clause[7][188] 	= partial_clause_prev[7][188] & 1'b1;
			partial_clause[7][189] 	= partial_clause_prev[7][189] & 1'b1;
			partial_clause[7][190] 	= partial_clause_prev[7][190] & 1'b1;
			partial_clause[7][191] 	= partial_clause_prev[7][191] & 1'b1;
			partial_clause[7][192] 	= partial_clause_prev[7][192] & 1'b1;
			partial_clause[7][193] 	= partial_clause_prev[7][193] & 1'b1;
			partial_clause[7][194] 	= partial_clause_prev[7][194] & 1'b1;
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & 1'b1;
			partial_clause[7][197] 	= partial_clause_prev[7][197] & 1'b1;
			partial_clause[7][198] 	= partial_clause_prev[7][198] & 1'b1;
			partial_clause[7][199] 	= partial_clause_prev[7][199] & x[54];
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & ~x[39] & ~x[40];
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & x[3];
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & x[57] & ~x[59];
			partial_clause[8][14] 	= partial_clause_prev[8][14] & x[32];
			partial_clause[8][15] 	= partial_clause_prev[8][15] & x[1];
			partial_clause[8][16] 	= partial_clause_prev[8][16] & x[2] & ~x[32];
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & x[4] & ~x[56];
			partial_clause[8][26] 	= partial_clause_prev[8][26] & x[3];
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & x[0] & ~x[30];
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & x[58] & ~x[61];
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & x[2];
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & ~x[1] & x[4];
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & ~x[13] & ~x[51];
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & x[3] & ~x[11];
			partial_clause[8][47] 	= partial_clause_prev[8][47] & x[33];
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & x[55];
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & ~x[29] & x[32];
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & x[31];
			partial_clause[8][70] 	= partial_clause_prev[8][70] & ~x[31];
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & x[3] & ~x[11] & ~x[40];
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & ~x[4];
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & x[4];
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & x[3] & ~x[14];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & x[2] & ~x[60];
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & x[1];
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			partial_clause[8][100] 	= partial_clause_prev[8][100] & 1'b1;
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & 1'b1;
			partial_clause[8][103] 	= partial_clause_prev[8][103] & 1'b1;
			partial_clause[8][104] 	= partial_clause_prev[8][104] & 1'b1;
			partial_clause[8][105] 	= partial_clause_prev[8][105] & x[23];
			partial_clause[8][106] 	= partial_clause_prev[8][106] & 1'b1;
			partial_clause[8][107] 	= partial_clause_prev[8][107] & 1'b1;
			partial_clause[8][108] 	= partial_clause_prev[8][108] & 1'b1;
			partial_clause[8][109] 	= partial_clause_prev[8][109] & ~x[2] & ~x[3];
			partial_clause[8][110] 	= partial_clause_prev[8][110] & x[52];
			partial_clause[8][111] 	= partial_clause_prev[8][111] & 1'b1;
			partial_clause[8][112] 	= partial_clause_prev[8][112] & 1'b1;
			partial_clause[8][113] 	= partial_clause_prev[8][113] & 1'b1;
			partial_clause[8][114] 	= partial_clause_prev[8][114] & 1'b1;
			partial_clause[8][115] 	= partial_clause_prev[8][115] & 1'b1;
			partial_clause[8][116] 	= partial_clause_prev[8][116] & 1'b1;
			partial_clause[8][117] 	= partial_clause_prev[8][117] & 1'b1;
			partial_clause[8][118] 	= partial_clause_prev[8][118] & 1'b1;
			partial_clause[8][119] 	= partial_clause_prev[8][119] & ~x[1] & ~x[2] & ~x[31] & ~x[32] & ~x[49];
			partial_clause[8][120] 	= partial_clause_prev[8][120] & 1'b1;
			partial_clause[8][121] 	= partial_clause_prev[8][121] & 1'b1;
			partial_clause[8][122] 	= partial_clause_prev[8][122] & 1'b1;
			partial_clause[8][123] 	= partial_clause_prev[8][123] & 1'b1;
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & 1'b1;
			partial_clause[8][126] 	= partial_clause_prev[8][126] & x[9];
			partial_clause[8][127] 	= partial_clause_prev[8][127] & x[37] & x[63];
			partial_clause[8][128] 	= partial_clause_prev[8][128] & x[8];
			partial_clause[8][129] 	= partial_clause_prev[8][129] & 1'b1;
			partial_clause[8][130] 	= partial_clause_prev[8][130] & 1'b1;
			partial_clause[8][131] 	= partial_clause_prev[8][131] & 1'b1;
			partial_clause[8][132] 	= partial_clause_prev[8][132] & ~x[23] & ~x[29] & ~x[55];
			partial_clause[8][133] 	= partial_clause_prev[8][133] & 1'b1;
			partial_clause[8][134] 	= partial_clause_prev[8][134] & 1'b1;
			partial_clause[8][135] 	= partial_clause_prev[8][135] & 1'b1;
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & x[9];
			partial_clause[8][138] 	= partial_clause_prev[8][138] & 1'b1;
			partial_clause[8][139] 	= partial_clause_prev[8][139] & x[34] & ~x[56];
			partial_clause[8][140] 	= partial_clause_prev[8][140] & 1'b1;
			partial_clause[8][141] 	= partial_clause_prev[8][141] & ~x[49];
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & 1'b1;
			partial_clause[8][144] 	= partial_clause_prev[8][144] & 1'b1;
			partial_clause[8][145] 	= partial_clause_prev[8][145] & 1'b1;
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & 1'b1;
			partial_clause[8][148] 	= partial_clause_prev[8][148] & x[37];
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & 1'b1;
			partial_clause[8][151] 	= partial_clause_prev[8][151] & x[48];
			partial_clause[8][152] 	= partial_clause_prev[8][152] & ~x[1] & ~x[3] & ~x[4] & ~x[5];
			partial_clause[8][153] 	= partial_clause_prev[8][153] & 1'b1;
			partial_clause[8][154] 	= partial_clause_prev[8][154] & 1'b1;
			partial_clause[8][155] 	= partial_clause_prev[8][155] & 1'b1;
			partial_clause[8][156] 	= partial_clause_prev[8][156] & 1'b1;
			partial_clause[8][157] 	= partial_clause_prev[8][157] & 1'b1;
			partial_clause[8][158] 	= partial_clause_prev[8][158] & 1'b1;
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & 1'b1;
			partial_clause[8][161] 	= partial_clause_prev[8][161] & 1'b1;
			partial_clause[8][162] 	= partial_clause_prev[8][162] & 1'b1;
			partial_clause[8][163] 	= partial_clause_prev[8][163] & 1'b1;
			partial_clause[8][164] 	= partial_clause_prev[8][164] & 1'b1;
			partial_clause[8][165] 	= partial_clause_prev[8][165] & 1'b1;
			partial_clause[8][166] 	= partial_clause_prev[8][166] & ~x[5];
			partial_clause[8][167] 	= partial_clause_prev[8][167] & x[7];
			partial_clause[8][168] 	= partial_clause_prev[8][168] & 1'b1;
			partial_clause[8][169] 	= partial_clause_prev[8][169] & 1'b1;
			partial_clause[8][170] 	= partial_clause_prev[8][170] & 1'b1;
			partial_clause[8][171] 	= partial_clause_prev[8][171] & 1'b1;
			partial_clause[8][172] 	= partial_clause_prev[8][172] & 1'b1;
			partial_clause[8][173] 	= partial_clause_prev[8][173] & 1'b1;
			partial_clause[8][174] 	= partial_clause_prev[8][174] & 1'b1;
			partial_clause[8][175] 	= partial_clause_prev[8][175] & 1'b1;
			partial_clause[8][176] 	= partial_clause_prev[8][176] & 1'b1;
			partial_clause[8][177] 	= partial_clause_prev[8][177] & 1'b1;
			partial_clause[8][178] 	= partial_clause_prev[8][178] & 1'b1;
			partial_clause[8][179] 	= partial_clause_prev[8][179] & x[6] & x[33];
			partial_clause[8][180] 	= partial_clause_prev[8][180] & 1'b1;
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & 1'b1;
			partial_clause[8][183] 	= partial_clause_prev[8][183] & 1'b1;
			partial_clause[8][184] 	= partial_clause_prev[8][184] & 1'b1;
			partial_clause[8][185] 	= partial_clause_prev[8][185] & 1'b1;
			partial_clause[8][186] 	= partial_clause_prev[8][186] & ~x[4];
			partial_clause[8][187] 	= partial_clause_prev[8][187] & 1'b1;
			partial_clause[8][188] 	= partial_clause_prev[8][188] & 1'b1;
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & ~x[29];
			partial_clause[8][191] 	= partial_clause_prev[8][191] & 1'b1;
			partial_clause[8][192] 	= partial_clause_prev[8][192] & 1'b1;
			partial_clause[8][193] 	= partial_clause_prev[8][193] & 1'b1;
			partial_clause[8][194] 	= partial_clause_prev[8][194] & 1'b1;
			partial_clause[8][195] 	= partial_clause_prev[8][195] & x[39];
			partial_clause[8][196] 	= partial_clause_prev[8][196] & 1'b1;
			partial_clause[8][197] 	= partial_clause_prev[8][197] & 1'b1;
			partial_clause[8][198] 	= partial_clause_prev[8][198] & 1'b1;
			partial_clause[8][199] 	= partial_clause_prev[8][199] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & x[19];
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & ~x[11];
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & ~x[59];
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & ~x[26] & ~x[58];
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & ~x[24];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & x[48];
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & ~x[10];
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & ~x[10];
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & ~x[31] & ~x[38];
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & ~x[56];
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & ~x[28];
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & ~x[28];
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & ~x[60] & ~x[62];
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & ~x[1];
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
			partial_clause[9][100] 	= partial_clause_prev[9][100] & 1'b1;
			partial_clause[9][101] 	= partial_clause_prev[9][101] & 1'b1;
			partial_clause[9][102] 	= partial_clause_prev[9][102] & 1'b1;
			partial_clause[9][103] 	= partial_clause_prev[9][103] & 1'b1;
			partial_clause[9][104] 	= partial_clause_prev[9][104] & 1'b1;
			partial_clause[9][105] 	= partial_clause_prev[9][105] & 1'b1;
			partial_clause[9][106] 	= partial_clause_prev[9][106] & 1'b1;
			partial_clause[9][107] 	= partial_clause_prev[9][107] & 1'b1;
			partial_clause[9][108] 	= partial_clause_prev[9][108] & 1'b1;
			partial_clause[9][109] 	= partial_clause_prev[9][109] & 1'b1;
			partial_clause[9][110] 	= partial_clause_prev[9][110] & x[42];
			partial_clause[9][111] 	= partial_clause_prev[9][111] & 1'b1;
			partial_clause[9][112] 	= partial_clause_prev[9][112] & 1'b1;
			partial_clause[9][113] 	= partial_clause_prev[9][113] & 1'b1;
			partial_clause[9][114] 	= partial_clause_prev[9][114] & 1'b1;
			partial_clause[9][115] 	= partial_clause_prev[9][115] & 1'b1;
			partial_clause[9][116] 	= partial_clause_prev[9][116] & 1'b1;
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & 1'b1;
			partial_clause[9][119] 	= partial_clause_prev[9][119] & 1'b1;
			partial_clause[9][120] 	= partial_clause_prev[9][120] & 1'b1;
			partial_clause[9][121] 	= partial_clause_prev[9][121] & 1'b1;
			partial_clause[9][122] 	= partial_clause_prev[9][122] & 1'b1;
			partial_clause[9][123] 	= partial_clause_prev[9][123] & 1'b1;
			partial_clause[9][124] 	= partial_clause_prev[9][124] & x[59];
			partial_clause[9][125] 	= partial_clause_prev[9][125] & 1'b1;
			partial_clause[9][126] 	= partial_clause_prev[9][126] & 1'b1;
			partial_clause[9][127] 	= partial_clause_prev[9][127] & 1'b1;
			partial_clause[9][128] 	= partial_clause_prev[9][128] & 1'b1;
			partial_clause[9][129] 	= partial_clause_prev[9][129] & ~x[2];
			partial_clause[9][130] 	= partial_clause_prev[9][130] & 1'b1;
			partial_clause[9][131] 	= partial_clause_prev[9][131] & 1'b1;
			partial_clause[9][132] 	= partial_clause_prev[9][132] & 1'b1;
			partial_clause[9][133] 	= partial_clause_prev[9][133] & x[58];
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & 1'b1;
			partial_clause[9][138] 	= partial_clause_prev[9][138] & 1'b1;
			partial_clause[9][139] 	= partial_clause_prev[9][139] & 1'b1;
			partial_clause[9][140] 	= partial_clause_prev[9][140] & 1'b1;
			partial_clause[9][141] 	= partial_clause_prev[9][141] & 1'b1;
			partial_clause[9][142] 	= partial_clause_prev[9][142] & 1'b1;
			partial_clause[9][143] 	= partial_clause_prev[9][143] & 1'b1;
			partial_clause[9][144] 	= partial_clause_prev[9][144] & 1'b1;
			partial_clause[9][145] 	= partial_clause_prev[9][145] & 1'b1;
			partial_clause[9][146] 	= partial_clause_prev[9][146] & 1'b1;
			partial_clause[9][147] 	= partial_clause_prev[9][147] & 1'b1;
			partial_clause[9][148] 	= partial_clause_prev[9][148] & 1'b1;
			partial_clause[9][149] 	= partial_clause_prev[9][149] & ~x[19];
			partial_clause[9][150] 	= partial_clause_prev[9][150] & 1'b1;
			partial_clause[9][151] 	= partial_clause_prev[9][151] & 1'b1;
			partial_clause[9][152] 	= partial_clause_prev[9][152] & 1'b1;
			partial_clause[9][153] 	= partial_clause_prev[9][153] & x[57];
			partial_clause[9][154] 	= partial_clause_prev[9][154] & 1'b1;
			partial_clause[9][155] 	= partial_clause_prev[9][155] & 1'b1;
			partial_clause[9][156] 	= partial_clause_prev[9][156] & 1'b1;
			partial_clause[9][157] 	= partial_clause_prev[9][157] & 1'b1;
			partial_clause[9][158] 	= partial_clause_prev[9][158] & 1'b1;
			partial_clause[9][159] 	= partial_clause_prev[9][159] & 1'b1;
			partial_clause[9][160] 	= partial_clause_prev[9][160] & 1'b1;
			partial_clause[9][161] 	= partial_clause_prev[9][161] & 1'b1;
			partial_clause[9][162] 	= partial_clause_prev[9][162] & 1'b1;
			partial_clause[9][163] 	= partial_clause_prev[9][163] & 1'b1;
			partial_clause[9][164] 	= partial_clause_prev[9][164] & 1'b1;
			partial_clause[9][165] 	= partial_clause_prev[9][165] & 1'b1;
			partial_clause[9][166] 	= partial_clause_prev[9][166] & 1'b1;
			partial_clause[9][167] 	= partial_clause_prev[9][167] & 1'b1;
			partial_clause[9][168] 	= partial_clause_prev[9][168] & 1'b1;
			partial_clause[9][169] 	= partial_clause_prev[9][169] & 1'b1;
			partial_clause[9][170] 	= partial_clause_prev[9][170] & 1'b1;
			partial_clause[9][171] 	= partial_clause_prev[9][171] & 1'b1;
			partial_clause[9][172] 	= partial_clause_prev[9][172] & 1'b1;
			partial_clause[9][173] 	= partial_clause_prev[9][173] & 1'b1;
			partial_clause[9][174] 	= partial_clause_prev[9][174] & 1'b1;
			partial_clause[9][175] 	= partial_clause_prev[9][175] & 1'b1;
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & x[57];
			partial_clause[9][178] 	= partial_clause_prev[9][178] & 1'b1;
			partial_clause[9][179] 	= partial_clause_prev[9][179] & x[57];
			partial_clause[9][180] 	= partial_clause_prev[9][180] & x[56];
			partial_clause[9][181] 	= partial_clause_prev[9][181] & 1'b1;
			partial_clause[9][182] 	= partial_clause_prev[9][182] & ~x[0];
			partial_clause[9][183] 	= partial_clause_prev[9][183] & 1'b1;
			partial_clause[9][184] 	= partial_clause_prev[9][184] & 1'b1;
			partial_clause[9][185] 	= partial_clause_prev[9][185] & 1'b1;
			partial_clause[9][186] 	= partial_clause_prev[9][186] & 1'b1;
			partial_clause[9][187] 	= partial_clause_prev[9][187] & 1'b1;
			partial_clause[9][188] 	= partial_clause_prev[9][188] & 1'b1;
			partial_clause[9][189] 	= partial_clause_prev[9][189] & x[2];
			partial_clause[9][190] 	= partial_clause_prev[9][190] & 1'b1;
			partial_clause[9][191] 	= partial_clause_prev[9][191] & 1'b1;
			partial_clause[9][192] 	= partial_clause_prev[9][192] & 1'b1;
			partial_clause[9][193] 	= partial_clause_prev[9][193] & 1'b1;
			partial_clause[9][194] 	= partial_clause_prev[9][194] & 1'b1;
			partial_clause[9][195] 	= partial_clause_prev[9][195] & x[60];
			partial_clause[9][196] 	= partial_clause_prev[9][196] & 1'b1;
			partial_clause[9][197] 	= partial_clause_prev[9][197] & 1'b1;
			partial_clause[9][198] 	= partial_clause_prev[9][198] & x[55];
			partial_clause[9][199] 	= partial_clause_prev[9][199] & 1'b1;
		end
	end
endmodule


module HCB_9 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & ~x[29];
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & x[53];
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & ~x[58];
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & ~x[32] & x[50];
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & ~x[3];
			partial_clause[0][28] 	= partial_clause_prev[0][28] & x[53];
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & x[49];
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & x[51];
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & x[51];
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & x[53];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & x[37];
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & ~x[19];
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			partial_clause[0][100] 	= partial_clause_prev[0][100] & 1'b1;
			partial_clause[0][101] 	= partial_clause_prev[0][101] & 1'b1;
			partial_clause[0][102] 	= partial_clause_prev[0][102] & ~x[43];
			partial_clause[0][103] 	= partial_clause_prev[0][103] & 1'b1;
			partial_clause[0][104] 	= partial_clause_prev[0][104] & 1'b1;
			partial_clause[0][105] 	= partial_clause_prev[0][105] & 1'b1;
			partial_clause[0][106] 	= partial_clause_prev[0][106] & x[7];
			partial_clause[0][107] 	= partial_clause_prev[0][107] & 1'b1;
			partial_clause[0][108] 	= partial_clause_prev[0][108] & ~x[19];
			partial_clause[0][109] 	= partial_clause_prev[0][109] & 1'b1;
			partial_clause[0][110] 	= partial_clause_prev[0][110] & 1'b1;
			partial_clause[0][111] 	= partial_clause_prev[0][111] & 1'b1;
			partial_clause[0][112] 	= partial_clause_prev[0][112] & 1'b1;
			partial_clause[0][113] 	= partial_clause_prev[0][113] & 1'b1;
			partial_clause[0][114] 	= partial_clause_prev[0][114] & 1'b1;
			partial_clause[0][115] 	= partial_clause_prev[0][115] & 1'b1;
			partial_clause[0][116] 	= partial_clause_prev[0][116] & 1'b1;
			partial_clause[0][117] 	= partial_clause_prev[0][117] & 1'b1;
			partial_clause[0][118] 	= partial_clause_prev[0][118] & 1'b1;
			partial_clause[0][119] 	= partial_clause_prev[0][119] & ~x[51];
			partial_clause[0][120] 	= partial_clause_prev[0][120] & 1'b1;
			partial_clause[0][121] 	= partial_clause_prev[0][121] & 1'b1;
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & 1'b1;
			partial_clause[0][124] 	= partial_clause_prev[0][124] & 1'b1;
			partial_clause[0][125] 	= partial_clause_prev[0][125] & 1'b1;
			partial_clause[0][126] 	= partial_clause_prev[0][126] & 1'b1;
			partial_clause[0][127] 	= partial_clause_prev[0][127] & 1'b1;
			partial_clause[0][128] 	= partial_clause_prev[0][128] & 1'b1;
			partial_clause[0][129] 	= partial_clause_prev[0][129] & 1'b1;
			partial_clause[0][130] 	= partial_clause_prev[0][130] & 1'b1;
			partial_clause[0][131] 	= partial_clause_prev[0][131] & 1'b1;
			partial_clause[0][132] 	= partial_clause_prev[0][132] & 1'b1;
			partial_clause[0][133] 	= partial_clause_prev[0][133] & 1'b1;
			partial_clause[0][134] 	= partial_clause_prev[0][134] & 1'b1;
			partial_clause[0][135] 	= partial_clause_prev[0][135] & 1'b1;
			partial_clause[0][136] 	= partial_clause_prev[0][136] & 1'b1;
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & 1'b1;
			partial_clause[0][139] 	= partial_clause_prev[0][139] & 1'b1;
			partial_clause[0][140] 	= partial_clause_prev[0][140] & 1'b1;
			partial_clause[0][141] 	= partial_clause_prev[0][141] & 1'b1;
			partial_clause[0][142] 	= partial_clause_prev[0][142] & 1'b1;
			partial_clause[0][143] 	= partial_clause_prev[0][143] & 1'b1;
			partial_clause[0][144] 	= partial_clause_prev[0][144] & 1'b1;
			partial_clause[0][145] 	= partial_clause_prev[0][145] & 1'b1;
			partial_clause[0][146] 	= partial_clause_prev[0][146] & 1'b1;
			partial_clause[0][147] 	= partial_clause_prev[0][147] & ~x[53];
			partial_clause[0][148] 	= partial_clause_prev[0][148] & 1'b1;
			partial_clause[0][149] 	= partial_clause_prev[0][149] & ~x[51] & ~x[53];
			partial_clause[0][150] 	= partial_clause_prev[0][150] & 1'b1;
			partial_clause[0][151] 	= partial_clause_prev[0][151] & x[60];
			partial_clause[0][152] 	= partial_clause_prev[0][152] & 1'b1;
			partial_clause[0][153] 	= partial_clause_prev[0][153] & 1'b1;
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & 1'b1;
			partial_clause[0][156] 	= partial_clause_prev[0][156] & 1'b1;
			partial_clause[0][157] 	= partial_clause_prev[0][157] & 1'b1;
			partial_clause[0][158] 	= partial_clause_prev[0][158] & 1'b1;
			partial_clause[0][159] 	= partial_clause_prev[0][159] & 1'b1;
			partial_clause[0][160] 	= partial_clause_prev[0][160] & 1'b1;
			partial_clause[0][161] 	= partial_clause_prev[0][161] & 1'b1;
			partial_clause[0][162] 	= partial_clause_prev[0][162] & 1'b1;
			partial_clause[0][163] 	= partial_clause_prev[0][163] & ~x[22];
			partial_clause[0][164] 	= partial_clause_prev[0][164] & 1'b1;
			partial_clause[0][165] 	= partial_clause_prev[0][165] & ~x[24];
			partial_clause[0][166] 	= partial_clause_prev[0][166] & 1'b1;
			partial_clause[0][167] 	= partial_clause_prev[0][167] & 1'b1;
			partial_clause[0][168] 	= partial_clause_prev[0][168] & 1'b1;
			partial_clause[0][169] 	= partial_clause_prev[0][169] & 1'b1;
			partial_clause[0][170] 	= partial_clause_prev[0][170] & 1'b1;
			partial_clause[0][171] 	= partial_clause_prev[0][171] & 1'b1;
			partial_clause[0][172] 	= partial_clause_prev[0][172] & x[33];
			partial_clause[0][173] 	= partial_clause_prev[0][173] & 1'b1;
			partial_clause[0][174] 	= partial_clause_prev[0][174] & 1'b1;
			partial_clause[0][175] 	= partial_clause_prev[0][175] & 1'b1;
			partial_clause[0][176] 	= partial_clause_prev[0][176] & 1'b1;
			partial_clause[0][177] 	= partial_clause_prev[0][177] & 1'b1;
			partial_clause[0][178] 	= partial_clause_prev[0][178] & 1'b1;
			partial_clause[0][179] 	= partial_clause_prev[0][179] & ~x[22];
			partial_clause[0][180] 	= partial_clause_prev[0][180] & 1'b1;
			partial_clause[0][181] 	= partial_clause_prev[0][181] & 1'b1;
			partial_clause[0][182] 	= partial_clause_prev[0][182] & 1'b1;
			partial_clause[0][183] 	= partial_clause_prev[0][183] & 1'b1;
			partial_clause[0][184] 	= partial_clause_prev[0][184] & 1'b1;
			partial_clause[0][185] 	= partial_clause_prev[0][185] & 1'b1;
			partial_clause[0][186] 	= partial_clause_prev[0][186] & 1'b1;
			partial_clause[0][187] 	= partial_clause_prev[0][187] & 1'b1;
			partial_clause[0][188] 	= partial_clause_prev[0][188] & 1'b1;
			partial_clause[0][189] 	= partial_clause_prev[0][189] & 1'b1;
			partial_clause[0][190] 	= partial_clause_prev[0][190] & 1'b1;
			partial_clause[0][191] 	= partial_clause_prev[0][191] & 1'b1;
			partial_clause[0][192] 	= partial_clause_prev[0][192] & 1'b1;
			partial_clause[0][193] 	= partial_clause_prev[0][193] & 1'b1;
			partial_clause[0][194] 	= partial_clause_prev[0][194] & 1'b1;
			partial_clause[0][195] 	= partial_clause_prev[0][195] & 1'b1;
			partial_clause[0][196] 	= partial_clause_prev[0][196] & ~x[5];
			partial_clause[0][197] 	= partial_clause_prev[0][197] & 1'b1;
			partial_clause[0][198] 	= partial_clause_prev[0][198] & 1'b1;
			partial_clause[0][199] 	= partial_clause_prev[0][199] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[2];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & ~x[27];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & ~x[21];
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & x[45];
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & x[41];
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & ~x[1];
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & x[10];
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & ~x[53];
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & x[14];
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & x[49];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & ~x[4] & ~x[53];
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & ~x[20];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & ~x[25] & ~x[27];
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & ~x[28];
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & x[45];
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & ~x[0];
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & x[42];
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			partial_clause[1][100] 	= partial_clause_prev[1][100] & 1'b1;
			partial_clause[1][101] 	= partial_clause_prev[1][101] & 1'b1;
			partial_clause[1][102] 	= partial_clause_prev[1][102] & ~x[32] & ~x[58];
			partial_clause[1][103] 	= partial_clause_prev[1][103] & 1'b1;
			partial_clause[1][104] 	= partial_clause_prev[1][104] & 1'b1;
			partial_clause[1][105] 	= partial_clause_prev[1][105] & 1'b1;
			partial_clause[1][106] 	= partial_clause_prev[1][106] & 1'b1;
			partial_clause[1][107] 	= partial_clause_prev[1][107] & ~x[48];
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & 1'b1;
			partial_clause[1][110] 	= partial_clause_prev[1][110] & ~x[2] & ~x[57] & ~x[58];
			partial_clause[1][111] 	= partial_clause_prev[1][111] & 1'b1;
			partial_clause[1][112] 	= partial_clause_prev[1][112] & ~x[58];
			partial_clause[1][113] 	= partial_clause_prev[1][113] & 1'b1;
			partial_clause[1][114] 	= partial_clause_prev[1][114] & 1'b1;
			partial_clause[1][115] 	= partial_clause_prev[1][115] & 1'b1;
			partial_clause[1][116] 	= partial_clause_prev[1][116] & x[0];
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & 1'b1;
			partial_clause[1][119] 	= partial_clause_prev[1][119] & 1'b1;
			partial_clause[1][120] 	= partial_clause_prev[1][120] & ~x[57];
			partial_clause[1][121] 	= partial_clause_prev[1][121] & 1'b1;
			partial_clause[1][122] 	= partial_clause_prev[1][122] & ~x[2];
			partial_clause[1][123] 	= partial_clause_prev[1][123] & ~x[28];
			partial_clause[1][124] 	= partial_clause_prev[1][124] & 1'b1;
			partial_clause[1][125] 	= partial_clause_prev[1][125] & ~x[31];
			partial_clause[1][126] 	= partial_clause_prev[1][126] & 1'b1;
			partial_clause[1][127] 	= partial_clause_prev[1][127] & 1'b1;
			partial_clause[1][128] 	= partial_clause_prev[1][128] & 1'b1;
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & 1'b1;
			partial_clause[1][131] 	= partial_clause_prev[1][131] & 1'b1;
			partial_clause[1][132] 	= partial_clause_prev[1][132] & 1'b1;
			partial_clause[1][133] 	= partial_clause_prev[1][133] & 1'b1;
			partial_clause[1][134] 	= partial_clause_prev[1][134] & 1'b1;
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & 1'b1;
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & ~x[30];
			partial_clause[1][139] 	= partial_clause_prev[1][139] & 1'b1;
			partial_clause[1][140] 	= partial_clause_prev[1][140] & 1'b1;
			partial_clause[1][141] 	= partial_clause_prev[1][141] & 1'b1;
			partial_clause[1][142] 	= partial_clause_prev[1][142] & 1'b1;
			partial_clause[1][143] 	= partial_clause_prev[1][143] & 1'b1;
			partial_clause[1][144] 	= partial_clause_prev[1][144] & 1'b1;
			partial_clause[1][145] 	= partial_clause_prev[1][145] & 1'b1;
			partial_clause[1][146] 	= partial_clause_prev[1][146] & 1'b1;
			partial_clause[1][147] 	= partial_clause_prev[1][147] & 1'b1;
			partial_clause[1][148] 	= partial_clause_prev[1][148] & 1'b1;
			partial_clause[1][149] 	= partial_clause_prev[1][149] & 1'b1;
			partial_clause[1][150] 	= partial_clause_prev[1][150] & ~x[9] & ~x[32];
			partial_clause[1][151] 	= partial_clause_prev[1][151] & 1'b1;
			partial_clause[1][152] 	= partial_clause_prev[1][152] & 1'b1;
			partial_clause[1][153] 	= partial_clause_prev[1][153] & 1'b1;
			partial_clause[1][154] 	= partial_clause_prev[1][154] & 1'b1;
			partial_clause[1][155] 	= partial_clause_prev[1][155] & x[53];
			partial_clause[1][156] 	= partial_clause_prev[1][156] & 1'b1;
			partial_clause[1][157] 	= partial_clause_prev[1][157] & 1'b1;
			partial_clause[1][158] 	= partial_clause_prev[1][158] & 1'b1;
			partial_clause[1][159] 	= partial_clause_prev[1][159] & ~x[3];
			partial_clause[1][160] 	= partial_clause_prev[1][160] & x[52];
			partial_clause[1][161] 	= partial_clause_prev[1][161] & 1'b1;
			partial_clause[1][162] 	= partial_clause_prev[1][162] & 1'b1;
			partial_clause[1][163] 	= partial_clause_prev[1][163] & ~x[30];
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & 1'b1;
			partial_clause[1][166] 	= partial_clause_prev[1][166] & 1'b1;
			partial_clause[1][167] 	= partial_clause_prev[1][167] & 1'b1;
			partial_clause[1][168] 	= partial_clause_prev[1][168] & x[24];
			partial_clause[1][169] 	= partial_clause_prev[1][169] & 1'b1;
			partial_clause[1][170] 	= partial_clause_prev[1][170] & 1'b1;
			partial_clause[1][171] 	= partial_clause_prev[1][171] & 1'b1;
			partial_clause[1][172] 	= partial_clause_prev[1][172] & 1'b1;
			partial_clause[1][173] 	= partial_clause_prev[1][173] & 1'b1;
			partial_clause[1][174] 	= partial_clause_prev[1][174] & 1'b1;
			partial_clause[1][175] 	= partial_clause_prev[1][175] & 1'b1;
			partial_clause[1][176] 	= partial_clause_prev[1][176] & 1'b1;
			partial_clause[1][177] 	= partial_clause_prev[1][177] & 1'b1;
			partial_clause[1][178] 	= partial_clause_prev[1][178] & 1'b1;
			partial_clause[1][179] 	= partial_clause_prev[1][179] & 1'b1;
			partial_clause[1][180] 	= partial_clause_prev[1][180] & 1'b1;
			partial_clause[1][181] 	= partial_clause_prev[1][181] & 1'b1;
			partial_clause[1][182] 	= partial_clause_prev[1][182] & 1'b1;
			partial_clause[1][183] 	= partial_clause_prev[1][183] & 1'b1;
			partial_clause[1][184] 	= partial_clause_prev[1][184] & 1'b1;
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & 1'b1;
			partial_clause[1][187] 	= partial_clause_prev[1][187] & 1'b1;
			partial_clause[1][188] 	= partial_clause_prev[1][188] & 1'b1;
			partial_clause[1][189] 	= partial_clause_prev[1][189] & 1'b1;
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & 1'b1;
			partial_clause[1][192] 	= partial_clause_prev[1][192] & 1'b1;
			partial_clause[1][193] 	= partial_clause_prev[1][193] & 1'b1;
			partial_clause[1][194] 	= partial_clause_prev[1][194] & 1'b1;
			partial_clause[1][195] 	= partial_clause_prev[1][195] & 1'b1;
			partial_clause[1][196] 	= partial_clause_prev[1][196] & 1'b1;
			partial_clause[1][197] 	= partial_clause_prev[1][197] & 1'b1;
			partial_clause[1][198] 	= partial_clause_prev[1][198] & 1'b1;
			partial_clause[1][199] 	= partial_clause_prev[1][199] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & ~x[54];
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & x[60];
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & ~x[25] & ~x[51] & ~x[56];
			partial_clause[2][17] 	= partial_clause_prev[2][17] & x[20];
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & x[36];
			partial_clause[2][20] 	= partial_clause_prev[2][20] & x[7];
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & ~x[31];
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & x[62];
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & x[4];
			partial_clause[2][41] 	= partial_clause_prev[2][41] & ~x[30] & ~x[56];
			partial_clause[2][42] 	= partial_clause_prev[2][42] & x[4];
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & x[30];
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & x[41];
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & x[35];
			partial_clause[2][61] 	= partial_clause_prev[2][61] & x[21];
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & ~x[55];
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & ~x[55];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & x[8];
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & x[34];
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & x[28];
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & x[32];
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & ~x[28] & ~x[57];
			partial_clause[2][99] 	= partial_clause_prev[2][99] & x[35];
			partial_clause[2][100] 	= partial_clause_prev[2][100] & ~x[33];
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & 1'b1;
			partial_clause[2][103] 	= partial_clause_prev[2][103] & 1'b1;
			partial_clause[2][104] 	= partial_clause_prev[2][104] & ~x[1] & ~x[3];
			partial_clause[2][105] 	= partial_clause_prev[2][105] & ~x[4];
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & 1'b1;
			partial_clause[2][108] 	= partial_clause_prev[2][108] & 1'b1;
			partial_clause[2][109] 	= partial_clause_prev[2][109] & 1'b1;
			partial_clause[2][110] 	= partial_clause_prev[2][110] & 1'b1;
			partial_clause[2][111] 	= partial_clause_prev[2][111] & 1'b1;
			partial_clause[2][112] 	= partial_clause_prev[2][112] & 1'b1;
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & 1'b1;
			partial_clause[2][115] 	= partial_clause_prev[2][115] & 1'b1;
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & 1'b1;
			partial_clause[2][118] 	= partial_clause_prev[2][118] & ~x[2] & ~x[3] & ~x[57];
			partial_clause[2][119] 	= partial_clause_prev[2][119] & 1'b1;
			partial_clause[2][120] 	= partial_clause_prev[2][120] & 1'b1;
			partial_clause[2][121] 	= partial_clause_prev[2][121] & 1'b1;
			partial_clause[2][122] 	= partial_clause_prev[2][122] & 1'b1;
			partial_clause[2][123] 	= partial_clause_prev[2][123] & 1'b1;
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & 1'b1;
			partial_clause[2][126] 	= partial_clause_prev[2][126] & 1'b1;
			partial_clause[2][127] 	= partial_clause_prev[2][127] & 1'b1;
			partial_clause[2][128] 	= partial_clause_prev[2][128] & 1'b1;
			partial_clause[2][129] 	= partial_clause_prev[2][129] & 1'b1;
			partial_clause[2][130] 	= partial_clause_prev[2][130] & 1'b1;
			partial_clause[2][131] 	= partial_clause_prev[2][131] & ~x[5];
			partial_clause[2][132] 	= partial_clause_prev[2][132] & 1'b1;
			partial_clause[2][133] 	= partial_clause_prev[2][133] & 1'b1;
			partial_clause[2][134] 	= partial_clause_prev[2][134] & 1'b1;
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & 1'b1;
			partial_clause[2][137] 	= partial_clause_prev[2][137] & 1'b1;
			partial_clause[2][138] 	= partial_clause_prev[2][138] & 1'b1;
			partial_clause[2][139] 	= partial_clause_prev[2][139] & 1'b1;
			partial_clause[2][140] 	= partial_clause_prev[2][140] & 1'b1;
			partial_clause[2][141] 	= partial_clause_prev[2][141] & ~x[33];
			partial_clause[2][142] 	= partial_clause_prev[2][142] & 1'b1;
			partial_clause[2][143] 	= partial_clause_prev[2][143] & 1'b1;
			partial_clause[2][144] 	= partial_clause_prev[2][144] & 1'b1;
			partial_clause[2][145] 	= partial_clause_prev[2][145] & 1'b1;
			partial_clause[2][146] 	= partial_clause_prev[2][146] & 1'b1;
			partial_clause[2][147] 	= partial_clause_prev[2][147] & 1'b1;
			partial_clause[2][148] 	= partial_clause_prev[2][148] & 1'b1;
			partial_clause[2][149] 	= partial_clause_prev[2][149] & 1'b1;
			partial_clause[2][150] 	= partial_clause_prev[2][150] & 1'b1;
			partial_clause[2][151] 	= partial_clause_prev[2][151] & 1'b1;
			partial_clause[2][152] 	= partial_clause_prev[2][152] & 1'b1;
			partial_clause[2][153] 	= partial_clause_prev[2][153] & 1'b1;
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & 1'b1;
			partial_clause[2][156] 	= partial_clause_prev[2][156] & 1'b1;
			partial_clause[2][157] 	= partial_clause_prev[2][157] & 1'b1;
			partial_clause[2][158] 	= partial_clause_prev[2][158] & 1'b1;
			partial_clause[2][159] 	= partial_clause_prev[2][159] & 1'b1;
			partial_clause[2][160] 	= partial_clause_prev[2][160] & 1'b1;
			partial_clause[2][161] 	= partial_clause_prev[2][161] & 1'b1;
			partial_clause[2][162] 	= partial_clause_prev[2][162] & ~x[4] & ~x[32];
			partial_clause[2][163] 	= partial_clause_prev[2][163] & 1'b1;
			partial_clause[2][164] 	= partial_clause_prev[2][164] & 1'b1;
			partial_clause[2][165] 	= partial_clause_prev[2][165] & 1'b1;
			partial_clause[2][166] 	= partial_clause_prev[2][166] & 1'b1;
			partial_clause[2][167] 	= partial_clause_prev[2][167] & 1'b1;
			partial_clause[2][168] 	= partial_clause_prev[2][168] & 1'b1;
			partial_clause[2][169] 	= partial_clause_prev[2][169] & ~x[3] & ~x[30] & ~x[58];
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & 1'b1;
			partial_clause[2][173] 	= partial_clause_prev[2][173] & 1'b1;
			partial_clause[2][174] 	= partial_clause_prev[2][174] & 1'b1;
			partial_clause[2][175] 	= partial_clause_prev[2][175] & 1'b1;
			partial_clause[2][176] 	= partial_clause_prev[2][176] & ~x[33];
			partial_clause[2][177] 	= partial_clause_prev[2][177] & 1'b1;
			partial_clause[2][178] 	= partial_clause_prev[2][178] & ~x[5];
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & 1'b1;
			partial_clause[2][181] 	= partial_clause_prev[2][181] & ~x[31];
			partial_clause[2][182] 	= partial_clause_prev[2][182] & 1'b1;
			partial_clause[2][183] 	= partial_clause_prev[2][183] & 1'b1;
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & 1'b1;
			partial_clause[2][186] 	= partial_clause_prev[2][186] & ~x[3];
			partial_clause[2][187] 	= partial_clause_prev[2][187] & 1'b1;
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & 1'b1;
			partial_clause[2][190] 	= partial_clause_prev[2][190] & 1'b1;
			partial_clause[2][191] 	= partial_clause_prev[2][191] & 1'b1;
			partial_clause[2][192] 	= partial_clause_prev[2][192] & 1'b1;
			partial_clause[2][193] 	= partial_clause_prev[2][193] & 1'b1;
			partial_clause[2][194] 	= partial_clause_prev[2][194] & 1'b1;
			partial_clause[2][195] 	= partial_clause_prev[2][195] & 1'b1;
			partial_clause[2][196] 	= partial_clause_prev[2][196] & 1'b1;
			partial_clause[2][197] 	= partial_clause_prev[2][197] & 1'b1;
			partial_clause[2][198] 	= partial_clause_prev[2][198] & ~x[2] & ~x[31] & ~x[57];
			partial_clause[2][199] 	= partial_clause_prev[2][199] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & x[26] & ~x[35] & x[51];
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & x[3] & x[57];
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & x[50];
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & x[56];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & ~x[6];
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & x[44];
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			partial_clause[3][100] 	= partial_clause_prev[3][100] & ~x[16];
			partial_clause[3][101] 	= partial_clause_prev[3][101] & 1'b1;
			partial_clause[3][102] 	= partial_clause_prev[3][102] & 1'b1;
			partial_clause[3][103] 	= partial_clause_prev[3][103] & 1'b1;
			partial_clause[3][104] 	= partial_clause_prev[3][104] & 1'b1;
			partial_clause[3][105] 	= partial_clause_prev[3][105] & 1'b1;
			partial_clause[3][106] 	= partial_clause_prev[3][106] & 1'b1;
			partial_clause[3][107] 	= partial_clause_prev[3][107] & 1'b1;
			partial_clause[3][108] 	= partial_clause_prev[3][108] & 1'b1;
			partial_clause[3][109] 	= partial_clause_prev[3][109] & 1'b1;
			partial_clause[3][110] 	= partial_clause_prev[3][110] & 1'b1;
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & 1'b1;
			partial_clause[3][113] 	= partial_clause_prev[3][113] & ~x[22];
			partial_clause[3][114] 	= partial_clause_prev[3][114] & 1'b1;
			partial_clause[3][115] 	= partial_clause_prev[3][115] & 1'b1;
			partial_clause[3][116] 	= partial_clause_prev[3][116] & 1'b1;
			partial_clause[3][117] 	= partial_clause_prev[3][117] & 1'b1;
			partial_clause[3][118] 	= partial_clause_prev[3][118] & 1'b1;
			partial_clause[3][119] 	= partial_clause_prev[3][119] & 1'b1;
			partial_clause[3][120] 	= partial_clause_prev[3][120] & 1'b1;
			partial_clause[3][121] 	= partial_clause_prev[3][121] & 1'b1;
			partial_clause[3][122] 	= partial_clause_prev[3][122] & 1'b1;
			partial_clause[3][123] 	= partial_clause_prev[3][123] & 1'b1;
			partial_clause[3][124] 	= partial_clause_prev[3][124] & 1'b1;
			partial_clause[3][125] 	= partial_clause_prev[3][125] & 1'b1;
			partial_clause[3][126] 	= partial_clause_prev[3][126] & 1'b1;
			partial_clause[3][127] 	= partial_clause_prev[3][127] & 1'b1;
			partial_clause[3][128] 	= partial_clause_prev[3][128] & 1'b1;
			partial_clause[3][129] 	= partial_clause_prev[3][129] & 1'b1;
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & 1'b1;
			partial_clause[3][132] 	= partial_clause_prev[3][132] & 1'b1;
			partial_clause[3][133] 	= partial_clause_prev[3][133] & 1'b1;
			partial_clause[3][134] 	= partial_clause_prev[3][134] & 1'b1;
			partial_clause[3][135] 	= partial_clause_prev[3][135] & 1'b1;
			partial_clause[3][136] 	= partial_clause_prev[3][136] & 1'b1;
			partial_clause[3][137] 	= partial_clause_prev[3][137] & 1'b1;
			partial_clause[3][138] 	= partial_clause_prev[3][138] & ~x[57];
			partial_clause[3][139] 	= partial_clause_prev[3][139] & ~x[49];
			partial_clause[3][140] 	= partial_clause_prev[3][140] & 1'b1;
			partial_clause[3][141] 	= partial_clause_prev[3][141] & x[62];
			partial_clause[3][142] 	= partial_clause_prev[3][142] & 1'b1;
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & ~x[20];
			partial_clause[3][145] 	= partial_clause_prev[3][145] & 1'b1;
			partial_clause[3][146] 	= partial_clause_prev[3][146] & 1'b1;
			partial_clause[3][147] 	= partial_clause_prev[3][147] & 1'b1;
			partial_clause[3][148] 	= partial_clause_prev[3][148] & 1'b1;
			partial_clause[3][149] 	= partial_clause_prev[3][149] & 1'b1;
			partial_clause[3][150] 	= partial_clause_prev[3][150] & 1'b1;
			partial_clause[3][151] 	= partial_clause_prev[3][151] & 1'b1;
			partial_clause[3][152] 	= partial_clause_prev[3][152] & 1'b1;
			partial_clause[3][153] 	= partial_clause_prev[3][153] & 1'b1;
			partial_clause[3][154] 	= partial_clause_prev[3][154] & 1'b1;
			partial_clause[3][155] 	= partial_clause_prev[3][155] & 1'b1;
			partial_clause[3][156] 	= partial_clause_prev[3][156] & ~x[1] & ~x[46];
			partial_clause[3][157] 	= partial_clause_prev[3][157] & 1'b1;
			partial_clause[3][158] 	= partial_clause_prev[3][158] & 1'b1;
			partial_clause[3][159] 	= partial_clause_prev[3][159] & 1'b1;
			partial_clause[3][160] 	= partial_clause_prev[3][160] & 1'b1;
			partial_clause[3][161] 	= partial_clause_prev[3][161] & 1'b1;
			partial_clause[3][162] 	= partial_clause_prev[3][162] & 1'b1;
			partial_clause[3][163] 	= partial_clause_prev[3][163] & x[8];
			partial_clause[3][164] 	= partial_clause_prev[3][164] & 1'b1;
			partial_clause[3][165] 	= partial_clause_prev[3][165] & 1'b1;
			partial_clause[3][166] 	= partial_clause_prev[3][166] & 1'b1;
			partial_clause[3][167] 	= partial_clause_prev[3][167] & 1'b1;
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & 1'b1;
			partial_clause[3][170] 	= partial_clause_prev[3][170] & 1'b1;
			partial_clause[3][171] 	= partial_clause_prev[3][171] & ~x[20];
			partial_clause[3][172] 	= partial_clause_prev[3][172] & 1'b1;
			partial_clause[3][173] 	= partial_clause_prev[3][173] & ~x[49];
			partial_clause[3][174] 	= partial_clause_prev[3][174] & 1'b1;
			partial_clause[3][175] 	= partial_clause_prev[3][175] & 1'b1;
			partial_clause[3][176] 	= partial_clause_prev[3][176] & 1'b1;
			partial_clause[3][177] 	= partial_clause_prev[3][177] & 1'b1;
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & 1'b1;
			partial_clause[3][180] 	= partial_clause_prev[3][180] & 1'b1;
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & 1'b1;
			partial_clause[3][183] 	= partial_clause_prev[3][183] & ~x[29] & ~x[57] & ~x[58];
			partial_clause[3][184] 	= partial_clause_prev[3][184] & 1'b1;
			partial_clause[3][185] 	= partial_clause_prev[3][185] & 1'b1;
			partial_clause[3][186] 	= partial_clause_prev[3][186] & 1'b1;
			partial_clause[3][187] 	= partial_clause_prev[3][187] & 1'b1;
			partial_clause[3][188] 	= partial_clause_prev[3][188] & 1'b1;
			partial_clause[3][189] 	= partial_clause_prev[3][189] & 1'b1;
			partial_clause[3][190] 	= partial_clause_prev[3][190] & 1'b1;
			partial_clause[3][191] 	= partial_clause_prev[3][191] & 1'b1;
			partial_clause[3][192] 	= partial_clause_prev[3][192] & 1'b1;
			partial_clause[3][193] 	= partial_clause_prev[3][193] & 1'b1;
			partial_clause[3][194] 	= partial_clause_prev[3][194] & 1'b1;
			partial_clause[3][195] 	= partial_clause_prev[3][195] & 1'b1;
			partial_clause[3][196] 	= partial_clause_prev[3][196] & 1'b1;
			partial_clause[3][197] 	= partial_clause_prev[3][197] & 1'b1;
			partial_clause[3][198] 	= partial_clause_prev[3][198] & 1'b1;
			partial_clause[3][199] 	= partial_clause_prev[3][199] & ~x[30];
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & x[35];
			partial_clause[4][2] 	= partial_clause_prev[4][2] & ~x[22];
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & ~x[24] & ~x[51];
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & ~x[52];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & 1'b1;
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & 1'b1;
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & ~x[51];
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & ~x[22];
			partial_clause[4][56] 	= partial_clause_prev[4][56] & x[14];
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & ~x[18] & ~x[26] & ~x[54];
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & x[10];
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			partial_clause[4][100] 	= partial_clause_prev[4][100] & 1'b1;
			partial_clause[4][101] 	= partial_clause_prev[4][101] & 1'b1;
			partial_clause[4][102] 	= partial_clause_prev[4][102] & 1'b1;
			partial_clause[4][103] 	= partial_clause_prev[4][103] & 1'b1;
			partial_clause[4][104] 	= partial_clause_prev[4][104] & x[24];
			partial_clause[4][105] 	= partial_clause_prev[4][105] & 1'b1;
			partial_clause[4][106] 	= partial_clause_prev[4][106] & 1'b1;
			partial_clause[4][107] 	= partial_clause_prev[4][107] & 1'b1;
			partial_clause[4][108] 	= partial_clause_prev[4][108] & 1'b1;
			partial_clause[4][109] 	= partial_clause_prev[4][109] & 1'b1;
			partial_clause[4][110] 	= partial_clause_prev[4][110] & 1'b1;
			partial_clause[4][111] 	= partial_clause_prev[4][111] & x[48];
			partial_clause[4][112] 	= partial_clause_prev[4][112] & 1'b1;
			partial_clause[4][113] 	= partial_clause_prev[4][113] & 1'b1;
			partial_clause[4][114] 	= partial_clause_prev[4][114] & x[17];
			partial_clause[4][115] 	= partial_clause_prev[4][115] & 1'b1;
			partial_clause[4][116] 	= partial_clause_prev[4][116] & 1'b1;
			partial_clause[4][117] 	= partial_clause_prev[4][117] & 1'b1;
			partial_clause[4][118] 	= partial_clause_prev[4][118] & 1'b1;
			partial_clause[4][119] 	= partial_clause_prev[4][119] & 1'b1;
			partial_clause[4][120] 	= partial_clause_prev[4][120] & 1'b1;
			partial_clause[4][121] 	= partial_clause_prev[4][121] & 1'b1;
			partial_clause[4][122] 	= partial_clause_prev[4][122] & 1'b1;
			partial_clause[4][123] 	= partial_clause_prev[4][123] & 1'b1;
			partial_clause[4][124] 	= partial_clause_prev[4][124] & 1'b1;
			partial_clause[4][125] 	= partial_clause_prev[4][125] & x[18];
			partial_clause[4][126] 	= partial_clause_prev[4][126] & 1'b1;
			partial_clause[4][127] 	= partial_clause_prev[4][127] & 1'b1;
			partial_clause[4][128] 	= partial_clause_prev[4][128] & 1'b1;
			partial_clause[4][129] 	= partial_clause_prev[4][129] & x[21];
			partial_clause[4][130] 	= partial_clause_prev[4][130] & 1'b1;
			partial_clause[4][131] 	= partial_clause_prev[4][131] & 1'b1;
			partial_clause[4][132] 	= partial_clause_prev[4][132] & 1'b1;
			partial_clause[4][133] 	= partial_clause_prev[4][133] & 1'b1;
			partial_clause[4][134] 	= partial_clause_prev[4][134] & 1'b1;
			partial_clause[4][135] 	= partial_clause_prev[4][135] & 1'b1;
			partial_clause[4][136] 	= partial_clause_prev[4][136] & x[19];
			partial_clause[4][137] 	= partial_clause_prev[4][137] & 1'b1;
			partial_clause[4][138] 	= partial_clause_prev[4][138] & 1'b1;
			partial_clause[4][139] 	= partial_clause_prev[4][139] & 1'b1;
			partial_clause[4][140] 	= partial_clause_prev[4][140] & x[25];
			partial_clause[4][141] 	= partial_clause_prev[4][141] & 1'b1;
			partial_clause[4][142] 	= partial_clause_prev[4][142] & x[19] & x[48];
			partial_clause[4][143] 	= partial_clause_prev[4][143] & 1'b1;
			partial_clause[4][144] 	= partial_clause_prev[4][144] & 1'b1;
			partial_clause[4][145] 	= partial_clause_prev[4][145] & 1'b1;
			partial_clause[4][146] 	= partial_clause_prev[4][146] & 1'b1;
			partial_clause[4][147] 	= partial_clause_prev[4][147] & 1'b1;
			partial_clause[4][148] 	= partial_clause_prev[4][148] & 1'b1;
			partial_clause[4][149] 	= partial_clause_prev[4][149] & 1'b1;
			partial_clause[4][150] 	= partial_clause_prev[4][150] & 1'b1;
			partial_clause[4][151] 	= partial_clause_prev[4][151] & 1'b1;
			partial_clause[4][152] 	= partial_clause_prev[4][152] & 1'b1;
			partial_clause[4][153] 	= partial_clause_prev[4][153] & 1'b1;
			partial_clause[4][154] 	= partial_clause_prev[4][154] & 1'b1;
			partial_clause[4][155] 	= partial_clause_prev[4][155] & 1'b1;
			partial_clause[4][156] 	= partial_clause_prev[4][156] & 1'b1;
			partial_clause[4][157] 	= partial_clause_prev[4][157] & 1'b1;
			partial_clause[4][158] 	= partial_clause_prev[4][158] & x[20];
			partial_clause[4][159] 	= partial_clause_prev[4][159] & x[23];
			partial_clause[4][160] 	= partial_clause_prev[4][160] & 1'b1;
			partial_clause[4][161] 	= partial_clause_prev[4][161] & 1'b1;
			partial_clause[4][162] 	= partial_clause_prev[4][162] & 1'b1;
			partial_clause[4][163] 	= partial_clause_prev[4][163] & 1'b1;
			partial_clause[4][164] 	= partial_clause_prev[4][164] & 1'b1;
			partial_clause[4][165] 	= partial_clause_prev[4][165] & x[1];
			partial_clause[4][166] 	= partial_clause_prev[4][166] & x[22];
			partial_clause[4][167] 	= partial_clause_prev[4][167] & x[27];
			partial_clause[4][168] 	= partial_clause_prev[4][168] & 1'b1;
			partial_clause[4][169] 	= partial_clause_prev[4][169] & x[52];
			partial_clause[4][170] 	= partial_clause_prev[4][170] & 1'b1;
			partial_clause[4][171] 	= partial_clause_prev[4][171] & x[2];
			partial_clause[4][172] 	= partial_clause_prev[4][172] & 1'b1;
			partial_clause[4][173] 	= partial_clause_prev[4][173] & 1'b1;
			partial_clause[4][174] 	= partial_clause_prev[4][174] & 1'b1;
			partial_clause[4][175] 	= partial_clause_prev[4][175] & 1'b1;
			partial_clause[4][176] 	= partial_clause_prev[4][176] & 1'b1;
			partial_clause[4][177] 	= partial_clause_prev[4][177] & 1'b1;
			partial_clause[4][178] 	= partial_clause_prev[4][178] & x[47];
			partial_clause[4][179] 	= partial_clause_prev[4][179] & 1'b1;
			partial_clause[4][180] 	= partial_clause_prev[4][180] & 1'b1;
			partial_clause[4][181] 	= partial_clause_prev[4][181] & 1'b1;
			partial_clause[4][182] 	= partial_clause_prev[4][182] & 1'b1;
			partial_clause[4][183] 	= partial_clause_prev[4][183] & 1'b1;
			partial_clause[4][184] 	= partial_clause_prev[4][184] & x[47];
			partial_clause[4][185] 	= partial_clause_prev[4][185] & 1'b1;
			partial_clause[4][186] 	= partial_clause_prev[4][186] & 1'b1;
			partial_clause[4][187] 	= partial_clause_prev[4][187] & 1'b1;
			partial_clause[4][188] 	= partial_clause_prev[4][188] & 1'b1;
			partial_clause[4][189] 	= partial_clause_prev[4][189] & 1'b1;
			partial_clause[4][190] 	= partial_clause_prev[4][190] & 1'b1;
			partial_clause[4][191] 	= partial_clause_prev[4][191] & 1'b1;
			partial_clause[4][192] 	= partial_clause_prev[4][192] & 1'b1;
			partial_clause[4][193] 	= partial_clause_prev[4][193] & x[54];
			partial_clause[4][194] 	= partial_clause_prev[4][194] & 1'b1;
			partial_clause[4][195] 	= partial_clause_prev[4][195] & 1'b1;
			partial_clause[4][196] 	= partial_clause_prev[4][196] & x[47];
			partial_clause[4][197] 	= partial_clause_prev[4][197] & 1'b1;
			partial_clause[4][198] 	= partial_clause_prev[4][198] & 1'b1;
			partial_clause[4][199] 	= partial_clause_prev[4][199] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & x[34];
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & x[36];
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & x[20];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & x[33];
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & x[53];
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & x[7];
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & x[57];
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			partial_clause[5][100] 	= partial_clause_prev[5][100] & 1'b1;
			partial_clause[5][101] 	= partial_clause_prev[5][101] & 1'b1;
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & 1'b1;
			partial_clause[5][104] 	= partial_clause_prev[5][104] & 1'b1;
			partial_clause[5][105] 	= partial_clause_prev[5][105] & 1'b1;
			partial_clause[5][106] 	= partial_clause_prev[5][106] & 1'b1;
			partial_clause[5][107] 	= partial_clause_prev[5][107] & 1'b1;
			partial_clause[5][108] 	= partial_clause_prev[5][108] & 1'b1;
			partial_clause[5][109] 	= partial_clause_prev[5][109] & 1'b1;
			partial_clause[5][110] 	= partial_clause_prev[5][110] & 1'b1;
			partial_clause[5][111] 	= partial_clause_prev[5][111] & 1'b1;
			partial_clause[5][112] 	= partial_clause_prev[5][112] & 1'b1;
			partial_clause[5][113] 	= partial_clause_prev[5][113] & 1'b1;
			partial_clause[5][114] 	= partial_clause_prev[5][114] & 1'b1;
			partial_clause[5][115] 	= partial_clause_prev[5][115] & 1'b1;
			partial_clause[5][116] 	= partial_clause_prev[5][116] & 1'b1;
			partial_clause[5][117] 	= partial_clause_prev[5][117] & 1'b1;
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & 1'b1;
			partial_clause[5][120] 	= partial_clause_prev[5][120] & 1'b1;
			partial_clause[5][121] 	= partial_clause_prev[5][121] & 1'b1;
			partial_clause[5][122] 	= partial_clause_prev[5][122] & 1'b1;
			partial_clause[5][123] 	= partial_clause_prev[5][123] & 1'b1;
			partial_clause[5][124] 	= partial_clause_prev[5][124] & 1'b1;
			partial_clause[5][125] 	= partial_clause_prev[5][125] & ~x[40];
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & 1'b1;
			partial_clause[5][128] 	= partial_clause_prev[5][128] & 1'b1;
			partial_clause[5][129] 	= partial_clause_prev[5][129] & 1'b1;
			partial_clause[5][130] 	= partial_clause_prev[5][130] & 1'b1;
			partial_clause[5][131] 	= partial_clause_prev[5][131] & 1'b1;
			partial_clause[5][132] 	= partial_clause_prev[5][132] & ~x[32] & ~x[49];
			partial_clause[5][133] 	= partial_clause_prev[5][133] & 1'b1;
			partial_clause[5][134] 	= partial_clause_prev[5][134] & 1'b1;
			partial_clause[5][135] 	= partial_clause_prev[5][135] & 1'b1;
			partial_clause[5][136] 	= partial_clause_prev[5][136] & 1'b1;
			partial_clause[5][137] 	= partial_clause_prev[5][137] & 1'b1;
			partial_clause[5][138] 	= partial_clause_prev[5][138] & 1'b1;
			partial_clause[5][139] 	= partial_clause_prev[5][139] & 1'b1;
			partial_clause[5][140] 	= partial_clause_prev[5][140] & 1'b1;
			partial_clause[5][141] 	= partial_clause_prev[5][141] & 1'b1;
			partial_clause[5][142] 	= partial_clause_prev[5][142] & 1'b1;
			partial_clause[5][143] 	= partial_clause_prev[5][143] & 1'b1;
			partial_clause[5][144] 	= partial_clause_prev[5][144] & 1'b1;
			partial_clause[5][145] 	= partial_clause_prev[5][145] & 1'b1;
			partial_clause[5][146] 	= partial_clause_prev[5][146] & 1'b1;
			partial_clause[5][147] 	= partial_clause_prev[5][147] & 1'b1;
			partial_clause[5][148] 	= partial_clause_prev[5][148] & 1'b1;
			partial_clause[5][149] 	= partial_clause_prev[5][149] & 1'b1;
			partial_clause[5][150] 	= partial_clause_prev[5][150] & 1'b1;
			partial_clause[5][151] 	= partial_clause_prev[5][151] & 1'b1;
			partial_clause[5][152] 	= partial_clause_prev[5][152] & 1'b1;
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & 1'b1;
			partial_clause[5][155] 	= partial_clause_prev[5][155] & 1'b1;
			partial_clause[5][156] 	= partial_clause_prev[5][156] & 1'b1;
			partial_clause[5][157] 	= partial_clause_prev[5][157] & 1'b1;
			partial_clause[5][158] 	= partial_clause_prev[5][158] & 1'b1;
			partial_clause[5][159] 	= partial_clause_prev[5][159] & 1'b1;
			partial_clause[5][160] 	= partial_clause_prev[5][160] & 1'b1;
			partial_clause[5][161] 	= partial_clause_prev[5][161] & 1'b1;
			partial_clause[5][162] 	= partial_clause_prev[5][162] & 1'b1;
			partial_clause[5][163] 	= partial_clause_prev[5][163] & 1'b1;
			partial_clause[5][164] 	= partial_clause_prev[5][164] & 1'b1;
			partial_clause[5][165] 	= partial_clause_prev[5][165] & 1'b1;
			partial_clause[5][166] 	= partial_clause_prev[5][166] & 1'b1;
			partial_clause[5][167] 	= partial_clause_prev[5][167] & x[42];
			partial_clause[5][168] 	= partial_clause_prev[5][168] & 1'b1;
			partial_clause[5][169] 	= partial_clause_prev[5][169] & 1'b1;
			partial_clause[5][170] 	= partial_clause_prev[5][170] & 1'b1;
			partial_clause[5][171] 	= partial_clause_prev[5][171] & 1'b1;
			partial_clause[5][172] 	= partial_clause_prev[5][172] & 1'b1;
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & 1'b1;
			partial_clause[5][175] 	= partial_clause_prev[5][175] & 1'b1;
			partial_clause[5][176] 	= partial_clause_prev[5][176] & 1'b1;
			partial_clause[5][177] 	= partial_clause_prev[5][177] & 1'b1;
			partial_clause[5][178] 	= partial_clause_prev[5][178] & 1'b1;
			partial_clause[5][179] 	= partial_clause_prev[5][179] & 1'b1;
			partial_clause[5][180] 	= partial_clause_prev[5][180] & 1'b1;
			partial_clause[5][181] 	= partial_clause_prev[5][181] & 1'b1;
			partial_clause[5][182] 	= partial_clause_prev[5][182] & 1'b1;
			partial_clause[5][183] 	= partial_clause_prev[5][183] & 1'b1;
			partial_clause[5][184] 	= partial_clause_prev[5][184] & 1'b1;
			partial_clause[5][185] 	= partial_clause_prev[5][185] & 1'b1;
			partial_clause[5][186] 	= partial_clause_prev[5][186] & 1'b1;
			partial_clause[5][187] 	= partial_clause_prev[5][187] & ~x[3];
			partial_clause[5][188] 	= partial_clause_prev[5][188] & 1'b1;
			partial_clause[5][189] 	= partial_clause_prev[5][189] & 1'b1;
			partial_clause[5][190] 	= partial_clause_prev[5][190] & 1'b1;
			partial_clause[5][191] 	= partial_clause_prev[5][191] & 1'b1;
			partial_clause[5][192] 	= partial_clause_prev[5][192] & 1'b1;
			partial_clause[5][193] 	= partial_clause_prev[5][193] & 1'b1;
			partial_clause[5][194] 	= partial_clause_prev[5][194] & 1'b1;
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & 1'b1;
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & 1'b1;
			partial_clause[5][199] 	= partial_clause_prev[5][199] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & x[26];
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & x[25];
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & ~x[50];
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & x[24];
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & x[27] & ~x[60];
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & x[42];
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & ~x[20] & x[25] & ~x[49];
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & x[0];
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			partial_clause[6][100] 	= partial_clause_prev[6][100] & ~x[0] & ~x[27];
			partial_clause[6][101] 	= partial_clause_prev[6][101] & 1'b1;
			partial_clause[6][102] 	= partial_clause_prev[6][102] & 1'b1;
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & 1'b1;
			partial_clause[6][105] 	= partial_clause_prev[6][105] & 1'b1;
			partial_clause[6][106] 	= partial_clause_prev[6][106] & 1'b1;
			partial_clause[6][107] 	= partial_clause_prev[6][107] & 1'b1;
			partial_clause[6][108] 	= partial_clause_prev[6][108] & x[20];
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & 1'b1;
			partial_clause[6][111] 	= partial_clause_prev[6][111] & 1'b1;
			partial_clause[6][112] 	= partial_clause_prev[6][112] & 1'b1;
			partial_clause[6][113] 	= partial_clause_prev[6][113] & 1'b1;
			partial_clause[6][114] 	= partial_clause_prev[6][114] & 1'b1;
			partial_clause[6][115] 	= partial_clause_prev[6][115] & 1'b1;
			partial_clause[6][116] 	= partial_clause_prev[6][116] & ~x[24];
			partial_clause[6][117] 	= partial_clause_prev[6][117] & ~x[22];
			partial_clause[6][118] 	= partial_clause_prev[6][118] & 1'b1;
			partial_clause[6][119] 	= partial_clause_prev[6][119] & x[46];
			partial_clause[6][120] 	= partial_clause_prev[6][120] & 1'b1;
			partial_clause[6][121] 	= partial_clause_prev[6][121] & 1'b1;
			partial_clause[6][122] 	= partial_clause_prev[6][122] & 1'b1;
			partial_clause[6][123] 	= partial_clause_prev[6][123] & ~x[28];
			partial_clause[6][124] 	= partial_clause_prev[6][124] & 1'b1;
			partial_clause[6][125] 	= partial_clause_prev[6][125] & 1'b1;
			partial_clause[6][126] 	= partial_clause_prev[6][126] & 1'b1;
			partial_clause[6][127] 	= partial_clause_prev[6][127] & 1'b1;
			partial_clause[6][128] 	= partial_clause_prev[6][128] & 1'b1;
			partial_clause[6][129] 	= partial_clause_prev[6][129] & 1'b1;
			partial_clause[6][130] 	= partial_clause_prev[6][130] & 1'b1;
			partial_clause[6][131] 	= partial_clause_prev[6][131] & 1'b1;
			partial_clause[6][132] 	= partial_clause_prev[6][132] & 1'b1;
			partial_clause[6][133] 	= partial_clause_prev[6][133] & 1'b1;
			partial_clause[6][134] 	= partial_clause_prev[6][134] & 1'b1;
			partial_clause[6][135] 	= partial_clause_prev[6][135] & 1'b1;
			partial_clause[6][136] 	= partial_clause_prev[6][136] & 1'b1;
			partial_clause[6][137] 	= partial_clause_prev[6][137] & 1'b1;
			partial_clause[6][138] 	= partial_clause_prev[6][138] & 1'b1;
			partial_clause[6][139] 	= partial_clause_prev[6][139] & 1'b1;
			partial_clause[6][140] 	= partial_clause_prev[6][140] & 1'b1;
			partial_clause[6][141] 	= partial_clause_prev[6][141] & 1'b1;
			partial_clause[6][142] 	= partial_clause_prev[6][142] & 1'b1;
			partial_clause[6][143] 	= partial_clause_prev[6][143] & 1'b1;
			partial_clause[6][144] 	= partial_clause_prev[6][144] & x[33];
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & 1'b1;
			partial_clause[6][147] 	= partial_clause_prev[6][147] & 1'b1;
			partial_clause[6][148] 	= partial_clause_prev[6][148] & 1'b1;
			partial_clause[6][149] 	= partial_clause_prev[6][149] & 1'b1;
			partial_clause[6][150] 	= partial_clause_prev[6][150] & 1'b1;
			partial_clause[6][151] 	= partial_clause_prev[6][151] & 1'b1;
			partial_clause[6][152] 	= partial_clause_prev[6][152] & ~x[22];
			partial_clause[6][153] 	= partial_clause_prev[6][153] & 1'b1;
			partial_clause[6][154] 	= partial_clause_prev[6][154] & 1'b1;
			partial_clause[6][155] 	= partial_clause_prev[6][155] & 1'b1;
			partial_clause[6][156] 	= partial_clause_prev[6][156] & 1'b1;
			partial_clause[6][157] 	= partial_clause_prev[6][157] & 1'b1;
			partial_clause[6][158] 	= partial_clause_prev[6][158] & x[48];
			partial_clause[6][159] 	= partial_clause_prev[6][159] & 1'b1;
			partial_clause[6][160] 	= partial_clause_prev[6][160] & 1'b1;
			partial_clause[6][161] 	= partial_clause_prev[6][161] & 1'b1;
			partial_clause[6][162] 	= partial_clause_prev[6][162] & x[16];
			partial_clause[6][163] 	= partial_clause_prev[6][163] & ~x[24];
			partial_clause[6][164] 	= partial_clause_prev[6][164] & 1'b1;
			partial_clause[6][165] 	= partial_clause_prev[6][165] & 1'b1;
			partial_clause[6][166] 	= partial_clause_prev[6][166] & 1'b1;
			partial_clause[6][167] 	= partial_clause_prev[6][167] & 1'b1;
			partial_clause[6][168] 	= partial_clause_prev[6][168] & 1'b1;
			partial_clause[6][169] 	= partial_clause_prev[6][169] & 1'b1;
			partial_clause[6][170] 	= partial_clause_prev[6][170] & x[17];
			partial_clause[6][171] 	= partial_clause_prev[6][171] & 1'b1;
			partial_clause[6][172] 	= partial_clause_prev[6][172] & 1'b1;
			partial_clause[6][173] 	= partial_clause_prev[6][173] & x[18];
			partial_clause[6][174] 	= partial_clause_prev[6][174] & 1'b1;
			partial_clause[6][175] 	= partial_clause_prev[6][175] & 1'b1;
			partial_clause[6][176] 	= partial_clause_prev[6][176] & 1'b1;
			partial_clause[6][177] 	= partial_clause_prev[6][177] & 1'b1;
			partial_clause[6][178] 	= partial_clause_prev[6][178] & 1'b1;
			partial_clause[6][179] 	= partial_clause_prev[6][179] & 1'b1;
			partial_clause[6][180] 	= partial_clause_prev[6][180] & x[18];
			partial_clause[6][181] 	= partial_clause_prev[6][181] & ~x[53];
			partial_clause[6][182] 	= partial_clause_prev[6][182] & ~x[25];
			partial_clause[6][183] 	= partial_clause_prev[6][183] & 1'b1;
			partial_clause[6][184] 	= partial_clause_prev[6][184] & 1'b1;
			partial_clause[6][185] 	= partial_clause_prev[6][185] & 1'b1;
			partial_clause[6][186] 	= partial_clause_prev[6][186] & 1'b1;
			partial_clause[6][187] 	= partial_clause_prev[6][187] & 1'b1;
			partial_clause[6][188] 	= partial_clause_prev[6][188] & 1'b1;
			partial_clause[6][189] 	= partial_clause_prev[6][189] & 1'b1;
			partial_clause[6][190] 	= partial_clause_prev[6][190] & 1'b1;
			partial_clause[6][191] 	= partial_clause_prev[6][191] & 1'b1;
			partial_clause[6][192] 	= partial_clause_prev[6][192] & 1'b1;
			partial_clause[6][193] 	= partial_clause_prev[6][193] & 1'b1;
			partial_clause[6][194] 	= partial_clause_prev[6][194] & 1'b1;
			partial_clause[6][195] 	= partial_clause_prev[6][195] & 1'b1;
			partial_clause[6][196] 	= partial_clause_prev[6][196] & 1'b1;
			partial_clause[6][197] 	= partial_clause_prev[6][197] & 1'b1;
			partial_clause[6][198] 	= partial_clause_prev[6][198] & 1'b1;
			partial_clause[6][199] 	= partial_clause_prev[6][199] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & ~x[22];
			partial_clause[7][10] 	= partial_clause_prev[7][10] & ~x[29] & x[50];
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & x[25];
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & ~x[50];
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & ~x[30];
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & ~x[1];
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & ~x[29];
			partial_clause[7][63] 	= partial_clause_prev[7][63] & ~x[20];
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & ~x[50];
			partial_clause[7][76] 	= partial_clause_prev[7][76] & ~x[48];
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & ~x[3] & x[25];
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & ~x[31];
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & ~x[5];
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & ~x[30];
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & ~x[1];
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & ~x[49];
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			partial_clause[7][100] 	= partial_clause_prev[7][100] & 1'b1;
			partial_clause[7][101] 	= partial_clause_prev[7][101] & 1'b1;
			partial_clause[7][102] 	= partial_clause_prev[7][102] & 1'b1;
			partial_clause[7][103] 	= partial_clause_prev[7][103] & x[5];
			partial_clause[7][104] 	= partial_clause_prev[7][104] & 1'b1;
			partial_clause[7][105] 	= partial_clause_prev[7][105] & 1'b1;
			partial_clause[7][106] 	= partial_clause_prev[7][106] & 1'b1;
			partial_clause[7][107] 	= partial_clause_prev[7][107] & 1'b1;
			partial_clause[7][108] 	= partial_clause_prev[7][108] & 1'b1;
			partial_clause[7][109] 	= partial_clause_prev[7][109] & 1'b1;
			partial_clause[7][110] 	= partial_clause_prev[7][110] & 1'b1;
			partial_clause[7][111] 	= partial_clause_prev[7][111] & x[2];
			partial_clause[7][112] 	= partial_clause_prev[7][112] & 1'b1;
			partial_clause[7][113] 	= partial_clause_prev[7][113] & 1'b1;
			partial_clause[7][114] 	= partial_clause_prev[7][114] & x[2];
			partial_clause[7][115] 	= partial_clause_prev[7][115] & x[20];
			partial_clause[7][116] 	= partial_clause_prev[7][116] & 1'b1;
			partial_clause[7][117] 	= partial_clause_prev[7][117] & 1'b1;
			partial_clause[7][118] 	= partial_clause_prev[7][118] & 1'b1;
			partial_clause[7][119] 	= partial_clause_prev[7][119] & 1'b1;
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & 1'b1;
			partial_clause[7][123] 	= partial_clause_prev[7][123] & 1'b1;
			partial_clause[7][124] 	= partial_clause_prev[7][124] & 1'b1;
			partial_clause[7][125] 	= partial_clause_prev[7][125] & x[3];
			partial_clause[7][126] 	= partial_clause_prev[7][126] & x[21] & x[23];
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & 1'b1;
			partial_clause[7][129] 	= partial_clause_prev[7][129] & 1'b1;
			partial_clause[7][130] 	= partial_clause_prev[7][130] & 1'b1;
			partial_clause[7][131] 	= partial_clause_prev[7][131] & 1'b1;
			partial_clause[7][132] 	= partial_clause_prev[7][132] & 1'b1;
			partial_clause[7][133] 	= partial_clause_prev[7][133] & 1'b1;
			partial_clause[7][134] 	= partial_clause_prev[7][134] & 1'b1;
			partial_clause[7][135] 	= partial_clause_prev[7][135] & 1'b1;
			partial_clause[7][136] 	= partial_clause_prev[7][136] & 1'b1;
			partial_clause[7][137] 	= partial_clause_prev[7][137] & 1'b1;
			partial_clause[7][138] 	= partial_clause_prev[7][138] & 1'b1;
			partial_clause[7][139] 	= partial_clause_prev[7][139] & 1'b1;
			partial_clause[7][140] 	= partial_clause_prev[7][140] & 1'b1;
			partial_clause[7][141] 	= partial_clause_prev[7][141] & 1'b1;
			partial_clause[7][142] 	= partial_clause_prev[7][142] & 1'b1;
			partial_clause[7][143] 	= partial_clause_prev[7][143] & 1'b1;
			partial_clause[7][144] 	= partial_clause_prev[7][144] & 1'b1;
			partial_clause[7][145] 	= partial_clause_prev[7][145] & 1'b1;
			partial_clause[7][146] 	= partial_clause_prev[7][146] & 1'b1;
			partial_clause[7][147] 	= partial_clause_prev[7][147] & 1'b1;
			partial_clause[7][148] 	= partial_clause_prev[7][148] & 1'b1;
			partial_clause[7][149] 	= partial_clause_prev[7][149] & 1'b1;
			partial_clause[7][150] 	= partial_clause_prev[7][150] & 1'b1;
			partial_clause[7][151] 	= partial_clause_prev[7][151] & 1'b1;
			partial_clause[7][152] 	= partial_clause_prev[7][152] & x[6];
			partial_clause[7][153] 	= partial_clause_prev[7][153] & 1'b1;
			partial_clause[7][154] 	= partial_clause_prev[7][154] & 1'b1;
			partial_clause[7][155] 	= partial_clause_prev[7][155] & 1'b1;
			partial_clause[7][156] 	= partial_clause_prev[7][156] & 1'b1;
			partial_clause[7][157] 	= partial_clause_prev[7][157] & 1'b1;
			partial_clause[7][158] 	= partial_clause_prev[7][158] & x[56];
			partial_clause[7][159] 	= partial_clause_prev[7][159] & x[27];
			partial_clause[7][160] 	= partial_clause_prev[7][160] & x[21];
			partial_clause[7][161] 	= partial_clause_prev[7][161] & 1'b1;
			partial_clause[7][162] 	= partial_clause_prev[7][162] & x[4];
			partial_clause[7][163] 	= partial_clause_prev[7][163] & 1'b1;
			partial_clause[7][164] 	= partial_clause_prev[7][164] & x[4];
			partial_clause[7][165] 	= partial_clause_prev[7][165] & 1'b1;
			partial_clause[7][166] 	= partial_clause_prev[7][166] & 1'b1;
			partial_clause[7][167] 	= partial_clause_prev[7][167] & 1'b1;
			partial_clause[7][168] 	= partial_clause_prev[7][168] & 1'b1;
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & 1'b1;
			partial_clause[7][171] 	= partial_clause_prev[7][171] & 1'b1;
			partial_clause[7][172] 	= partial_clause_prev[7][172] & 1'b1;
			partial_clause[7][173] 	= partial_clause_prev[7][173] & 1'b1;
			partial_clause[7][174] 	= partial_clause_prev[7][174] & 1'b1;
			partial_clause[7][175] 	= partial_clause_prev[7][175] & 1'b1;
			partial_clause[7][176] 	= partial_clause_prev[7][176] & 1'b1;
			partial_clause[7][177] 	= partial_clause_prev[7][177] & 1'b1;
			partial_clause[7][178] 	= partial_clause_prev[7][178] & 1'b1;
			partial_clause[7][179] 	= partial_clause_prev[7][179] & 1'b1;
			partial_clause[7][180] 	= partial_clause_prev[7][180] & 1'b1;
			partial_clause[7][181] 	= partial_clause_prev[7][181] & 1'b1;
			partial_clause[7][182] 	= partial_clause_prev[7][182] & 1'b1;
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & 1'b1;
			partial_clause[7][185] 	= partial_clause_prev[7][185] & 1'b1;
			partial_clause[7][186] 	= partial_clause_prev[7][186] & 1'b1;
			partial_clause[7][187] 	= partial_clause_prev[7][187] & 1'b1;
			partial_clause[7][188] 	= partial_clause_prev[7][188] & 1'b1;
			partial_clause[7][189] 	= partial_clause_prev[7][189] & x[19];
			partial_clause[7][190] 	= partial_clause_prev[7][190] & 1'b1;
			partial_clause[7][191] 	= partial_clause_prev[7][191] & x[31];
			partial_clause[7][192] 	= partial_clause_prev[7][192] & 1'b1;
			partial_clause[7][193] 	= partial_clause_prev[7][193] & 1'b1;
			partial_clause[7][194] 	= partial_clause_prev[7][194] & 1'b1;
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & 1'b1;
			partial_clause[7][197] 	= partial_clause_prev[7][197] & 1'b1;
			partial_clause[7][198] 	= partial_clause_prev[7][198] & 1'b1;
			partial_clause[7][199] 	= partial_clause_prev[7][199] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & ~x[3];
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & ~x[21];
			partial_clause[8][6] 	= partial_clause_prev[8][6] & x[46];
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & ~x[20];
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & ~x[33];
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & x[11];
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & ~x[33];
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & x[12];
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & ~x[21];
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & ~x[61];
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & x[61];
			partial_clause[8][87] 	= partial_clause_prev[8][87] & ~x[61];
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & x[15];
			partial_clause[8][100] 	= partial_clause_prev[8][100] & 1'b1;
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & 1'b1;
			partial_clause[8][103] 	= partial_clause_prev[8][103] & 1'b1;
			partial_clause[8][104] 	= partial_clause_prev[8][104] & 1'b1;
			partial_clause[8][105] 	= partial_clause_prev[8][105] & 1'b1;
			partial_clause[8][106] 	= partial_clause_prev[8][106] & 1'b1;
			partial_clause[8][107] 	= partial_clause_prev[8][107] & 1'b1;
			partial_clause[8][108] 	= partial_clause_prev[8][108] & 1'b1;
			partial_clause[8][109] 	= partial_clause_prev[8][109] & 1'b1;
			partial_clause[8][110] 	= partial_clause_prev[8][110] & 1'b1;
			partial_clause[8][111] 	= partial_clause_prev[8][111] & 1'b1;
			partial_clause[8][112] 	= partial_clause_prev[8][112] & 1'b1;
			partial_clause[8][113] 	= partial_clause_prev[8][113] & ~x[52] & ~x[60];
			partial_clause[8][114] 	= partial_clause_prev[8][114] & ~x[32] & ~x[60];
			partial_clause[8][115] 	= partial_clause_prev[8][115] & 1'b1;
			partial_clause[8][116] 	= partial_clause_prev[8][116] & 1'b1;
			partial_clause[8][117] 	= partial_clause_prev[8][117] & x[63];
			partial_clause[8][118] 	= partial_clause_prev[8][118] & 1'b1;
			partial_clause[8][119] 	= partial_clause_prev[8][119] & 1'b1;
			partial_clause[8][120] 	= partial_clause_prev[8][120] & 1'b1;
			partial_clause[8][121] 	= partial_clause_prev[8][121] & 1'b1;
			partial_clause[8][122] 	= partial_clause_prev[8][122] & 1'b1;
			partial_clause[8][123] 	= partial_clause_prev[8][123] & 1'b1;
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & 1'b1;
			partial_clause[8][126] 	= partial_clause_prev[8][126] & 1'b1;
			partial_clause[8][127] 	= partial_clause_prev[8][127] & 1'b1;
			partial_clause[8][128] 	= partial_clause_prev[8][128] & 1'b1;
			partial_clause[8][129] 	= partial_clause_prev[8][129] & 1'b1;
			partial_clause[8][130] 	= partial_clause_prev[8][130] & 1'b1;
			partial_clause[8][131] 	= partial_clause_prev[8][131] & 1'b1;
			partial_clause[8][132] 	= partial_clause_prev[8][132] & 1'b1;
			partial_clause[8][133] 	= partial_clause_prev[8][133] & 1'b1;
			partial_clause[8][134] 	= partial_clause_prev[8][134] & 1'b1;
			partial_clause[8][135] 	= partial_clause_prev[8][135] & ~x[53] & ~x[61];
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & 1'b1;
			partial_clause[8][138] 	= partial_clause_prev[8][138] & 1'b1;
			partial_clause[8][139] 	= partial_clause_prev[8][139] & ~x[19] & ~x[30] & ~x[57] & ~x[58];
			partial_clause[8][140] 	= partial_clause_prev[8][140] & x[14];
			partial_clause[8][141] 	= partial_clause_prev[8][141] & ~x[53];
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & 1'b1;
			partial_clause[8][144] 	= partial_clause_prev[8][144] & 1'b1;
			partial_clause[8][145] 	= partial_clause_prev[8][145] & 1'b1;
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & 1'b1;
			partial_clause[8][148] 	= partial_clause_prev[8][148] & 1'b1;
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & 1'b1;
			partial_clause[8][151] 	= partial_clause_prev[8][151] & 1'b1;
			partial_clause[8][152] 	= partial_clause_prev[8][152] & 1'b1;
			partial_clause[8][153] 	= partial_clause_prev[8][153] & 1'b1;
			partial_clause[8][154] 	= partial_clause_prev[8][154] & 1'b1;
			partial_clause[8][155] 	= partial_clause_prev[8][155] & 1'b1;
			partial_clause[8][156] 	= partial_clause_prev[8][156] & 1'b1;
			partial_clause[8][157] 	= partial_clause_prev[8][157] & 1'b1;
			partial_clause[8][158] 	= partial_clause_prev[8][158] & 1'b1;
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & 1'b1;
			partial_clause[8][161] 	= partial_clause_prev[8][161] & 1'b1;
			partial_clause[8][162] 	= partial_clause_prev[8][162] & 1'b1;
			partial_clause[8][163] 	= partial_clause_prev[8][163] & 1'b1;
			partial_clause[8][164] 	= partial_clause_prev[8][164] & 1'b1;
			partial_clause[8][165] 	= partial_clause_prev[8][165] & ~x[52];
			partial_clause[8][166] 	= partial_clause_prev[8][166] & 1'b1;
			partial_clause[8][167] 	= partial_clause_prev[8][167] & ~x[30] & ~x[59];
			partial_clause[8][168] 	= partial_clause_prev[8][168] & 1'b1;
			partial_clause[8][169] 	= partial_clause_prev[8][169] & 1'b1;
			partial_clause[8][170] 	= partial_clause_prev[8][170] & 1'b1;
			partial_clause[8][171] 	= partial_clause_prev[8][171] & 1'b1;
			partial_clause[8][172] 	= partial_clause_prev[8][172] & 1'b1;
			partial_clause[8][173] 	= partial_clause_prev[8][173] & 1'b1;
			partial_clause[8][174] 	= partial_clause_prev[8][174] & 1'b1;
			partial_clause[8][175] 	= partial_clause_prev[8][175] & 1'b1;
			partial_clause[8][176] 	= partial_clause_prev[8][176] & 1'b1;
			partial_clause[8][177] 	= partial_clause_prev[8][177] & 1'b1;
			partial_clause[8][178] 	= partial_clause_prev[8][178] & 1'b1;
			partial_clause[8][179] 	= partial_clause_prev[8][179] & ~x[56];
			partial_clause[8][180] 	= partial_clause_prev[8][180] & 1'b1;
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & 1'b1;
			partial_clause[8][183] 	= partial_clause_prev[8][183] & 1'b1;
			partial_clause[8][184] 	= partial_clause_prev[8][184] & 1'b1;
			partial_clause[8][185] 	= partial_clause_prev[8][185] & 1'b1;
			partial_clause[8][186] 	= partial_clause_prev[8][186] & 1'b1;
			partial_clause[8][187] 	= partial_clause_prev[8][187] & 1'b1;
			partial_clause[8][188] 	= partial_clause_prev[8][188] & 1'b1;
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & ~x[33] & ~x[56];
			partial_clause[8][191] 	= partial_clause_prev[8][191] & 1'b1;
			partial_clause[8][192] 	= partial_clause_prev[8][192] & 1'b1;
			partial_clause[8][193] 	= partial_clause_prev[8][193] & 1'b1;
			partial_clause[8][194] 	= partial_clause_prev[8][194] & ~x[48] & ~x[50] & ~x[58];
			partial_clause[8][195] 	= partial_clause_prev[8][195] & 1'b1;
			partial_clause[8][196] 	= partial_clause_prev[8][196] & 1'b1;
			partial_clause[8][197] 	= partial_clause_prev[8][197] & x[36];
			partial_clause[8][198] 	= partial_clause_prev[8][198] & 1'b1;
			partial_clause[8][199] 	= partial_clause_prev[8][199] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & ~x[46];
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & ~x[3];
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & ~x[20] & ~x[22];
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & ~x[24];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & ~x[24] & ~x[51];
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & ~x[19];
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & x[10];
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & ~x[29];
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & ~x[23];
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & ~x[18];
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & ~x[23] & ~x[50];
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & x[15];
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
			partial_clause[9][100] 	= partial_clause_prev[9][100] & 1'b1;
			partial_clause[9][101] 	= partial_clause_prev[9][101] & 1'b1;
			partial_clause[9][102] 	= partial_clause_prev[9][102] & 1'b1;
			partial_clause[9][103] 	= partial_clause_prev[9][103] & 1'b1;
			partial_clause[9][104] 	= partial_clause_prev[9][104] & 1'b1;
			partial_clause[9][105] 	= partial_clause_prev[9][105] & 1'b1;
			partial_clause[9][106] 	= partial_clause_prev[9][106] & 1'b1;
			partial_clause[9][107] 	= partial_clause_prev[9][107] & 1'b1;
			partial_clause[9][108] 	= partial_clause_prev[9][108] & 1'b1;
			partial_clause[9][109] 	= partial_clause_prev[9][109] & 1'b1;
			partial_clause[9][110] 	= partial_clause_prev[9][110] & 1'b1;
			partial_clause[9][111] 	= partial_clause_prev[9][111] & 1'b1;
			partial_clause[9][112] 	= partial_clause_prev[9][112] & 1'b1;
			partial_clause[9][113] 	= partial_clause_prev[9][113] & 1'b1;
			partial_clause[9][114] 	= partial_clause_prev[9][114] & 1'b1;
			partial_clause[9][115] 	= partial_clause_prev[9][115] & 1'b1;
			partial_clause[9][116] 	= partial_clause_prev[9][116] & 1'b1;
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & ~x[62];
			partial_clause[9][119] 	= partial_clause_prev[9][119] & 1'b1;
			partial_clause[9][120] 	= partial_clause_prev[9][120] & 1'b1;
			partial_clause[9][121] 	= partial_clause_prev[9][121] & 1'b1;
			partial_clause[9][122] 	= partial_clause_prev[9][122] & 1'b1;
			partial_clause[9][123] 	= partial_clause_prev[9][123] & 1'b1;
			partial_clause[9][124] 	= partial_clause_prev[9][124] & 1'b1;
			partial_clause[9][125] 	= partial_clause_prev[9][125] & 1'b1;
			partial_clause[9][126] 	= partial_clause_prev[9][126] & 1'b1;
			partial_clause[9][127] 	= partial_clause_prev[9][127] & 1'b1;
			partial_clause[9][128] 	= partial_clause_prev[9][128] & 1'b1;
			partial_clause[9][129] 	= partial_clause_prev[9][129] & 1'b1;
			partial_clause[9][130] 	= partial_clause_prev[9][130] & 1'b1;
			partial_clause[9][131] 	= partial_clause_prev[9][131] & 1'b1;
			partial_clause[9][132] 	= partial_clause_prev[9][132] & 1'b1;
			partial_clause[9][133] 	= partial_clause_prev[9][133] & 1'b1;
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & 1'b1;
			partial_clause[9][138] 	= partial_clause_prev[9][138] & 1'b1;
			partial_clause[9][139] 	= partial_clause_prev[9][139] & x[19];
			partial_clause[9][140] 	= partial_clause_prev[9][140] & 1'b1;
			partial_clause[9][141] 	= partial_clause_prev[9][141] & x[20];
			partial_clause[9][142] 	= partial_clause_prev[9][142] & 1'b1;
			partial_clause[9][143] 	= partial_clause_prev[9][143] & 1'b1;
			partial_clause[9][144] 	= partial_clause_prev[9][144] & 1'b1;
			partial_clause[9][145] 	= partial_clause_prev[9][145] & 1'b1;
			partial_clause[9][146] 	= partial_clause_prev[9][146] & 1'b1;
			partial_clause[9][147] 	= partial_clause_prev[9][147] & 1'b1;
			partial_clause[9][148] 	= partial_clause_prev[9][148] & 1'b1;
			partial_clause[9][149] 	= partial_clause_prev[9][149] & 1'b1;
			partial_clause[9][150] 	= partial_clause_prev[9][150] & 1'b1;
			partial_clause[9][151] 	= partial_clause_prev[9][151] & 1'b1;
			partial_clause[9][152] 	= partial_clause_prev[9][152] & 1'b1;
			partial_clause[9][153] 	= partial_clause_prev[9][153] & 1'b1;
			partial_clause[9][154] 	= partial_clause_prev[9][154] & 1'b1;
			partial_clause[9][155] 	= partial_clause_prev[9][155] & 1'b1;
			partial_clause[9][156] 	= partial_clause_prev[9][156] & 1'b1;
			partial_clause[9][157] 	= partial_clause_prev[9][157] & 1'b1;
			partial_clause[9][158] 	= partial_clause_prev[9][158] & 1'b1;
			partial_clause[9][159] 	= partial_clause_prev[9][159] & 1'b1;
			partial_clause[9][160] 	= partial_clause_prev[9][160] & x[50];
			partial_clause[9][161] 	= partial_clause_prev[9][161] & 1'b1;
			partial_clause[9][162] 	= partial_clause_prev[9][162] & 1'b1;
			partial_clause[9][163] 	= partial_clause_prev[9][163] & 1'b1;
			partial_clause[9][164] 	= partial_clause_prev[9][164] & ~x[63];
			partial_clause[9][165] 	= partial_clause_prev[9][165] & 1'b1;
			partial_clause[9][166] 	= partial_clause_prev[9][166] & 1'b1;
			partial_clause[9][167] 	= partial_clause_prev[9][167] & 1'b1;
			partial_clause[9][168] 	= partial_clause_prev[9][168] & x[24];
			partial_clause[9][169] 	= partial_clause_prev[9][169] & 1'b1;
			partial_clause[9][170] 	= partial_clause_prev[9][170] & 1'b1;
			partial_clause[9][171] 	= partial_clause_prev[9][171] & x[18];
			partial_clause[9][172] 	= partial_clause_prev[9][172] & 1'b1;
			partial_clause[9][173] 	= partial_clause_prev[9][173] & 1'b1;
			partial_clause[9][174] 	= partial_clause_prev[9][174] & 1'b1;
			partial_clause[9][175] 	= partial_clause_prev[9][175] & 1'b1;
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & 1'b1;
			partial_clause[9][178] 	= partial_clause_prev[9][178] & 1'b1;
			partial_clause[9][179] 	= partial_clause_prev[9][179] & 1'b1;
			partial_clause[9][180] 	= partial_clause_prev[9][180] & 1'b1;
			partial_clause[9][181] 	= partial_clause_prev[9][181] & 1'b1;
			partial_clause[9][182] 	= partial_clause_prev[9][182] & 1'b1;
			partial_clause[9][183] 	= partial_clause_prev[9][183] & 1'b1;
			partial_clause[9][184] 	= partial_clause_prev[9][184] & 1'b1;
			partial_clause[9][185] 	= partial_clause_prev[9][185] & 1'b1;
			partial_clause[9][186] 	= partial_clause_prev[9][186] & 1'b1;
			partial_clause[9][187] 	= partial_clause_prev[9][187] & 1'b1;
			partial_clause[9][188] 	= partial_clause_prev[9][188] & x[55] & x[56];
			partial_clause[9][189] 	= partial_clause_prev[9][189] & 1'b1;
			partial_clause[9][190] 	= partial_clause_prev[9][190] & 1'b1;
			partial_clause[9][191] 	= partial_clause_prev[9][191] & 1'b1;
			partial_clause[9][192] 	= partial_clause_prev[9][192] & 1'b1;
			partial_clause[9][193] 	= partial_clause_prev[9][193] & 1'b1;
			partial_clause[9][194] 	= partial_clause_prev[9][194] & 1'b1;
			partial_clause[9][195] 	= partial_clause_prev[9][195] & 1'b1;
			partial_clause[9][196] 	= partial_clause_prev[9][196] & 1'b1;
			partial_clause[9][197] 	= partial_clause_prev[9][197] & 1'b1;
			partial_clause[9][198] 	= partial_clause_prev[9][198] & 1'b1;
			partial_clause[9][199] 	= partial_clause_prev[9][199] & 1'b1;
		end
	end
endmodule


module HCB_10 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & x[14];
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & x[16];
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & ~x[61];
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & x[15];
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			partial_clause[0][100] 	= partial_clause_prev[0][100] & 1'b1;
			partial_clause[0][101] 	= partial_clause_prev[0][101] & 1'b1;
			partial_clause[0][102] 	= partial_clause_prev[0][102] & 1'b1;
			partial_clause[0][103] 	= partial_clause_prev[0][103] & 1'b1;
			partial_clause[0][104] 	= partial_clause_prev[0][104] & 1'b1;
			partial_clause[0][105] 	= partial_clause_prev[0][105] & 1'b1;
			partial_clause[0][106] 	= partial_clause_prev[0][106] & 1'b1;
			partial_clause[0][107] 	= partial_clause_prev[0][107] & 1'b1;
			partial_clause[0][108] 	= partial_clause_prev[0][108] & 1'b1;
			partial_clause[0][109] 	= partial_clause_prev[0][109] & 1'b1;
			partial_clause[0][110] 	= partial_clause_prev[0][110] & 1'b1;
			partial_clause[0][111] 	= partial_clause_prev[0][111] & 1'b1;
			partial_clause[0][112] 	= partial_clause_prev[0][112] & 1'b1;
			partial_clause[0][113] 	= partial_clause_prev[0][113] & 1'b1;
			partial_clause[0][114] 	= partial_clause_prev[0][114] & 1'b1;
			partial_clause[0][115] 	= partial_clause_prev[0][115] & 1'b1;
			partial_clause[0][116] 	= partial_clause_prev[0][116] & 1'b1;
			partial_clause[0][117] 	= partial_clause_prev[0][117] & 1'b1;
			partial_clause[0][118] 	= partial_clause_prev[0][118] & x[51];
			partial_clause[0][119] 	= partial_clause_prev[0][119] & ~x[16];
			partial_clause[0][120] 	= partial_clause_prev[0][120] & 1'b1;
			partial_clause[0][121] 	= partial_clause_prev[0][121] & 1'b1;
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & 1'b1;
			partial_clause[0][124] 	= partial_clause_prev[0][124] & x[48];
			partial_clause[0][125] 	= partial_clause_prev[0][125] & ~x[7];
			partial_clause[0][126] 	= partial_clause_prev[0][126] & 1'b1;
			partial_clause[0][127] 	= partial_clause_prev[0][127] & 1'b1;
			partial_clause[0][128] 	= partial_clause_prev[0][128] & 1'b1;
			partial_clause[0][129] 	= partial_clause_prev[0][129] & 1'b1;
			partial_clause[0][130] 	= partial_clause_prev[0][130] & 1'b1;
			partial_clause[0][131] 	= partial_clause_prev[0][131] & 1'b1;
			partial_clause[0][132] 	= partial_clause_prev[0][132] & 1'b1;
			partial_clause[0][133] 	= partial_clause_prev[0][133] & 1'b1;
			partial_clause[0][134] 	= partial_clause_prev[0][134] & 1'b1;
			partial_clause[0][135] 	= partial_clause_prev[0][135] & 1'b1;
			partial_clause[0][136] 	= partial_clause_prev[0][136] & ~x[29];
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & 1'b1;
			partial_clause[0][139] 	= partial_clause_prev[0][139] & 1'b1;
			partial_clause[0][140] 	= partial_clause_prev[0][140] & 1'b1;
			partial_clause[0][141] 	= partial_clause_prev[0][141] & 1'b1;
			partial_clause[0][142] 	= partial_clause_prev[0][142] & 1'b1;
			partial_clause[0][143] 	= partial_clause_prev[0][143] & 1'b1;
			partial_clause[0][144] 	= partial_clause_prev[0][144] & 1'b1;
			partial_clause[0][145] 	= partial_clause_prev[0][145] & 1'b1;
			partial_clause[0][146] 	= partial_clause_prev[0][146] & 1'b1;
			partial_clause[0][147] 	= partial_clause_prev[0][147] & 1'b1;
			partial_clause[0][148] 	= partial_clause_prev[0][148] & 1'b1;
			partial_clause[0][149] 	= partial_clause_prev[0][149] & ~x[17];
			partial_clause[0][150] 	= partial_clause_prev[0][150] & 1'b1;
			partial_clause[0][151] 	= partial_clause_prev[0][151] & 1'b1;
			partial_clause[0][152] 	= partial_clause_prev[0][152] & 1'b1;
			partial_clause[0][153] 	= partial_clause_prev[0][153] & 1'b1;
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & 1'b1;
			partial_clause[0][156] 	= partial_clause_prev[0][156] & 1'b1;
			partial_clause[0][157] 	= partial_clause_prev[0][157] & ~x[17];
			partial_clause[0][158] 	= partial_clause_prev[0][158] & 1'b1;
			partial_clause[0][159] 	= partial_clause_prev[0][159] & 1'b1;
			partial_clause[0][160] 	= partial_clause_prev[0][160] & 1'b1;
			partial_clause[0][161] 	= partial_clause_prev[0][161] & ~x[44];
			partial_clause[0][162] 	= partial_clause_prev[0][162] & 1'b1;
			partial_clause[0][163] 	= partial_clause_prev[0][163] & 1'b1;
			partial_clause[0][164] 	= partial_clause_prev[0][164] & 1'b1;
			partial_clause[0][165] 	= partial_clause_prev[0][165] & 1'b1;
			partial_clause[0][166] 	= partial_clause_prev[0][166] & 1'b1;
			partial_clause[0][167] 	= partial_clause_prev[0][167] & ~x[6] & ~x[13] & ~x[18];
			partial_clause[0][168] 	= partial_clause_prev[0][168] & 1'b1;
			partial_clause[0][169] 	= partial_clause_prev[0][169] & 1'b1;
			partial_clause[0][170] 	= partial_clause_prev[0][170] & 1'b1;
			partial_clause[0][171] 	= partial_clause_prev[0][171] & 1'b1;
			partial_clause[0][172] 	= partial_clause_prev[0][172] & 1'b1;
			partial_clause[0][173] 	= partial_clause_prev[0][173] & ~x[17];
			partial_clause[0][174] 	= partial_clause_prev[0][174] & 1'b1;
			partial_clause[0][175] 	= partial_clause_prev[0][175] & 1'b1;
			partial_clause[0][176] 	= partial_clause_prev[0][176] & 1'b1;
			partial_clause[0][177] 	= partial_clause_prev[0][177] & 1'b1;
			partial_clause[0][178] 	= partial_clause_prev[0][178] & 1'b1;
			partial_clause[0][179] 	= partial_clause_prev[0][179] & 1'b1;
			partial_clause[0][180] 	= partial_clause_prev[0][180] & 1'b1;
			partial_clause[0][181] 	= partial_clause_prev[0][181] & 1'b1;
			partial_clause[0][182] 	= partial_clause_prev[0][182] & 1'b1;
			partial_clause[0][183] 	= partial_clause_prev[0][183] & 1'b1;
			partial_clause[0][184] 	= partial_clause_prev[0][184] & 1'b1;
			partial_clause[0][185] 	= partial_clause_prev[0][185] & 1'b1;
			partial_clause[0][186] 	= partial_clause_prev[0][186] & 1'b1;
			partial_clause[0][187] 	= partial_clause_prev[0][187] & 1'b1;
			partial_clause[0][188] 	= partial_clause_prev[0][188] & 1'b1;
			partial_clause[0][189] 	= partial_clause_prev[0][189] & 1'b1;
			partial_clause[0][190] 	= partial_clause_prev[0][190] & 1'b1;
			partial_clause[0][191] 	= partial_clause_prev[0][191] & 1'b1;
			partial_clause[0][192] 	= partial_clause_prev[0][192] & 1'b1;
			partial_clause[0][193] 	= partial_clause_prev[0][193] & 1'b1;
			partial_clause[0][194] 	= partial_clause_prev[0][194] & 1'b1;
			partial_clause[0][195] 	= partial_clause_prev[0][195] & 1'b1;
			partial_clause[0][196] 	= partial_clause_prev[0][196] & 1'b1;
			partial_clause[0][197] 	= partial_clause_prev[0][197] & 1'b1;
			partial_clause[0][198] 	= partial_clause_prev[0][198] & 1'b1;
			partial_clause[0][199] 	= partial_clause_prev[0][199] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & ~x[12];
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & x[60];
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & x[34];
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & x[1];
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & 1'b1;
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & ~x[53];
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & 1'b1;
			partial_clause[1][75] 	= partial_clause_prev[1][75] & x[60];
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & x[0];
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & ~x[44];
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			partial_clause[1][100] 	= partial_clause_prev[1][100] & 1'b1;
			partial_clause[1][101] 	= partial_clause_prev[1][101] & 1'b1;
			partial_clause[1][102] 	= partial_clause_prev[1][102] & 1'b1;
			partial_clause[1][103] 	= partial_clause_prev[1][103] & 1'b1;
			partial_clause[1][104] 	= partial_clause_prev[1][104] & 1'b1;
			partial_clause[1][105] 	= partial_clause_prev[1][105] & 1'b1;
			partial_clause[1][106] 	= partial_clause_prev[1][106] & 1'b1;
			partial_clause[1][107] 	= partial_clause_prev[1][107] & 1'b1;
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & 1'b1;
			partial_clause[1][110] 	= partial_clause_prev[1][110] & 1'b1;
			partial_clause[1][111] 	= partial_clause_prev[1][111] & x[16];
			partial_clause[1][112] 	= partial_clause_prev[1][112] & ~x[21];
			partial_clause[1][113] 	= partial_clause_prev[1][113] & 1'b1;
			partial_clause[1][114] 	= partial_clause_prev[1][114] & 1'b1;
			partial_clause[1][115] 	= partial_clause_prev[1][115] & 1'b1;
			partial_clause[1][116] 	= partial_clause_prev[1][116] & 1'b1;
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & 1'b1;
			partial_clause[1][119] 	= partial_clause_prev[1][119] & 1'b1;
			partial_clause[1][120] 	= partial_clause_prev[1][120] & ~x[21];
			partial_clause[1][121] 	= partial_clause_prev[1][121] & 1'b1;
			partial_clause[1][122] 	= partial_clause_prev[1][122] & 1'b1;
			partial_clause[1][123] 	= partial_clause_prev[1][123] & 1'b1;
			partial_clause[1][124] 	= partial_clause_prev[1][124] & 1'b1;
			partial_clause[1][125] 	= partial_clause_prev[1][125] & 1'b1;
			partial_clause[1][126] 	= partial_clause_prev[1][126] & 1'b1;
			partial_clause[1][127] 	= partial_clause_prev[1][127] & 1'b1;
			partial_clause[1][128] 	= partial_clause_prev[1][128] & ~x[8];
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & 1'b1;
			partial_clause[1][131] 	= partial_clause_prev[1][131] & 1'b1;
			partial_clause[1][132] 	= partial_clause_prev[1][132] & 1'b1;
			partial_clause[1][133] 	= partial_clause_prev[1][133] & 1'b1;
			partial_clause[1][134] 	= partial_clause_prev[1][134] & 1'b1;
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & 1'b1;
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & 1'b1;
			partial_clause[1][139] 	= partial_clause_prev[1][139] & 1'b1;
			partial_clause[1][140] 	= partial_clause_prev[1][140] & 1'b1;
			partial_clause[1][141] 	= partial_clause_prev[1][141] & 1'b1;
			partial_clause[1][142] 	= partial_clause_prev[1][142] & 1'b1;
			partial_clause[1][143] 	= partial_clause_prev[1][143] & 1'b1;
			partial_clause[1][144] 	= partial_clause_prev[1][144] & 1'b1;
			partial_clause[1][145] 	= partial_clause_prev[1][145] & 1'b1;
			partial_clause[1][146] 	= partial_clause_prev[1][146] & 1'b1;
			partial_clause[1][147] 	= partial_clause_prev[1][147] & 1'b1;
			partial_clause[1][148] 	= partial_clause_prev[1][148] & 1'b1;
			partial_clause[1][149] 	= partial_clause_prev[1][149] & 1'b1;
			partial_clause[1][150] 	= partial_clause_prev[1][150] & 1'b1;
			partial_clause[1][151] 	= partial_clause_prev[1][151] & 1'b1;
			partial_clause[1][152] 	= partial_clause_prev[1][152] & 1'b1;
			partial_clause[1][153] 	= partial_clause_prev[1][153] & 1'b1;
			partial_clause[1][154] 	= partial_clause_prev[1][154] & 1'b1;
			partial_clause[1][155] 	= partial_clause_prev[1][155] & 1'b1;
			partial_clause[1][156] 	= partial_clause_prev[1][156] & 1'b1;
			partial_clause[1][157] 	= partial_clause_prev[1][157] & 1'b1;
			partial_clause[1][158] 	= partial_clause_prev[1][158] & 1'b1;
			partial_clause[1][159] 	= partial_clause_prev[1][159] & 1'b1;
			partial_clause[1][160] 	= partial_clause_prev[1][160] & 1'b1;
			partial_clause[1][161] 	= partial_clause_prev[1][161] & 1'b1;
			partial_clause[1][162] 	= partial_clause_prev[1][162] & 1'b1;
			partial_clause[1][163] 	= partial_clause_prev[1][163] & 1'b1;
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & 1'b1;
			partial_clause[1][166] 	= partial_clause_prev[1][166] & 1'b1;
			partial_clause[1][167] 	= partial_clause_prev[1][167] & 1'b1;
			partial_clause[1][168] 	= partial_clause_prev[1][168] & 1'b1;
			partial_clause[1][169] 	= partial_clause_prev[1][169] & 1'b1;
			partial_clause[1][170] 	= partial_clause_prev[1][170] & 1'b1;
			partial_clause[1][171] 	= partial_clause_prev[1][171] & 1'b1;
			partial_clause[1][172] 	= partial_clause_prev[1][172] & 1'b1;
			partial_clause[1][173] 	= partial_clause_prev[1][173] & 1'b1;
			partial_clause[1][174] 	= partial_clause_prev[1][174] & 1'b1;
			partial_clause[1][175] 	= partial_clause_prev[1][175] & 1'b1;
			partial_clause[1][176] 	= partial_clause_prev[1][176] & 1'b1;
			partial_clause[1][177] 	= partial_clause_prev[1][177] & 1'b1;
			partial_clause[1][178] 	= partial_clause_prev[1][178] & 1'b1;
			partial_clause[1][179] 	= partial_clause_prev[1][179] & 1'b1;
			partial_clause[1][180] 	= partial_clause_prev[1][180] & 1'b1;
			partial_clause[1][181] 	= partial_clause_prev[1][181] & 1'b1;
			partial_clause[1][182] 	= partial_clause_prev[1][182] & 1'b1;
			partial_clause[1][183] 	= partial_clause_prev[1][183] & 1'b1;
			partial_clause[1][184] 	= partial_clause_prev[1][184] & 1'b1;
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & 1'b1;
			partial_clause[1][187] 	= partial_clause_prev[1][187] & 1'b1;
			partial_clause[1][188] 	= partial_clause_prev[1][188] & 1'b1;
			partial_clause[1][189] 	= partial_clause_prev[1][189] & 1'b1;
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & 1'b1;
			partial_clause[1][192] 	= partial_clause_prev[1][192] & 1'b1;
			partial_clause[1][193] 	= partial_clause_prev[1][193] & 1'b1;
			partial_clause[1][194] 	= partial_clause_prev[1][194] & 1'b1;
			partial_clause[1][195] 	= partial_clause_prev[1][195] & 1'b1;
			partial_clause[1][196] 	= partial_clause_prev[1][196] & 1'b1;
			partial_clause[1][197] 	= partial_clause_prev[1][197] & 1'b1;
			partial_clause[1][198] 	= partial_clause_prev[1][198] & 1'b1;
			partial_clause[1][199] 	= partial_clause_prev[1][199] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & x[58];
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & ~x[49];
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & x[25];
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & ~x[18];
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & x[57];
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & x[3];
			partial_clause[2][63] 	= partial_clause_prev[2][63] & ~x[49];
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & ~x[18] & ~x[48];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & x[26];
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & ~x[12];
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & x[0];
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			partial_clause[2][100] 	= partial_clause_prev[2][100] & 1'b1;
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & 1'b1;
			partial_clause[2][103] 	= partial_clause_prev[2][103] & 1'b1;
			partial_clause[2][104] 	= partial_clause_prev[2][104] & ~x[21];
			partial_clause[2][105] 	= partial_clause_prev[2][105] & 1'b1;
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & 1'b1;
			partial_clause[2][108] 	= partial_clause_prev[2][108] & 1'b1;
			partial_clause[2][109] 	= partial_clause_prev[2][109] & 1'b1;
			partial_clause[2][110] 	= partial_clause_prev[2][110] & 1'b1;
			partial_clause[2][111] 	= partial_clause_prev[2][111] & 1'b1;
			partial_clause[2][112] 	= partial_clause_prev[2][112] & 1'b1;
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & 1'b1;
			partial_clause[2][115] 	= partial_clause_prev[2][115] & 1'b1;
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & 1'b1;
			partial_clause[2][118] 	= partial_clause_prev[2][118] & 1'b1;
			partial_clause[2][119] 	= partial_clause_prev[2][119] & 1'b1;
			partial_clause[2][120] 	= partial_clause_prev[2][120] & 1'b1;
			partial_clause[2][121] 	= partial_clause_prev[2][121] & 1'b1;
			partial_clause[2][122] 	= partial_clause_prev[2][122] & 1'b1;
			partial_clause[2][123] 	= partial_clause_prev[2][123] & 1'b1;
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & 1'b1;
			partial_clause[2][126] 	= partial_clause_prev[2][126] & 1'b1;
			partial_clause[2][127] 	= partial_clause_prev[2][127] & 1'b1;
			partial_clause[2][128] 	= partial_clause_prev[2][128] & 1'b1;
			partial_clause[2][129] 	= partial_clause_prev[2][129] & 1'b1;
			partial_clause[2][130] 	= partial_clause_prev[2][130] & 1'b1;
			partial_clause[2][131] 	= partial_clause_prev[2][131] & ~x[24];
			partial_clause[2][132] 	= partial_clause_prev[2][132] & 1'b1;
			partial_clause[2][133] 	= partial_clause_prev[2][133] & 1'b1;
			partial_clause[2][134] 	= partial_clause_prev[2][134] & 1'b1;
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & x[44];
			partial_clause[2][137] 	= partial_clause_prev[2][137] & 1'b1;
			partial_clause[2][138] 	= partial_clause_prev[2][138] & 1'b1;
			partial_clause[2][139] 	= partial_clause_prev[2][139] & 1'b1;
			partial_clause[2][140] 	= partial_clause_prev[2][140] & 1'b1;
			partial_clause[2][141] 	= partial_clause_prev[2][141] & 1'b1;
			partial_clause[2][142] 	= partial_clause_prev[2][142] & 1'b1;
			partial_clause[2][143] 	= partial_clause_prev[2][143] & x[42];
			partial_clause[2][144] 	= partial_clause_prev[2][144] & 1'b1;
			partial_clause[2][145] 	= partial_clause_prev[2][145] & 1'b1;
			partial_clause[2][146] 	= partial_clause_prev[2][146] & 1'b1;
			partial_clause[2][147] 	= partial_clause_prev[2][147] & 1'b1;
			partial_clause[2][148] 	= partial_clause_prev[2][148] & 1'b1;
			partial_clause[2][149] 	= partial_clause_prev[2][149] & 1'b1;
			partial_clause[2][150] 	= partial_clause_prev[2][150] & 1'b1;
			partial_clause[2][151] 	= partial_clause_prev[2][151] & 1'b1;
			partial_clause[2][152] 	= partial_clause_prev[2][152] & 1'b1;
			partial_clause[2][153] 	= partial_clause_prev[2][153] & x[45];
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & 1'b1;
			partial_clause[2][156] 	= partial_clause_prev[2][156] & 1'b1;
			partial_clause[2][157] 	= partial_clause_prev[2][157] & 1'b1;
			partial_clause[2][158] 	= partial_clause_prev[2][158] & 1'b1;
			partial_clause[2][159] 	= partial_clause_prev[2][159] & 1'b1;
			partial_clause[2][160] 	= partial_clause_prev[2][160] & 1'b1;
			partial_clause[2][161] 	= partial_clause_prev[2][161] & ~x[49];
			partial_clause[2][162] 	= partial_clause_prev[2][162] & 1'b1;
			partial_clause[2][163] 	= partial_clause_prev[2][163] & x[47];
			partial_clause[2][164] 	= partial_clause_prev[2][164] & 1'b1;
			partial_clause[2][165] 	= partial_clause_prev[2][165] & 1'b1;
			partial_clause[2][166] 	= partial_clause_prev[2][166] & 1'b1;
			partial_clause[2][167] 	= partial_clause_prev[2][167] & 1'b1;
			partial_clause[2][168] 	= partial_clause_prev[2][168] & 1'b1;
			partial_clause[2][169] 	= partial_clause_prev[2][169] & 1'b1;
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & 1'b1;
			partial_clause[2][173] 	= partial_clause_prev[2][173] & 1'b1;
			partial_clause[2][174] 	= partial_clause_prev[2][174] & 1'b1;
			partial_clause[2][175] 	= partial_clause_prev[2][175] & 1'b1;
			partial_clause[2][176] 	= partial_clause_prev[2][176] & 1'b1;
			partial_clause[2][177] 	= partial_clause_prev[2][177] & x[15];
			partial_clause[2][178] 	= partial_clause_prev[2][178] & 1'b1;
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & 1'b1;
			partial_clause[2][181] 	= partial_clause_prev[2][181] & 1'b1;
			partial_clause[2][182] 	= partial_clause_prev[2][182] & 1'b1;
			partial_clause[2][183] 	= partial_clause_prev[2][183] & 1'b1;
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & 1'b1;
			partial_clause[2][186] 	= partial_clause_prev[2][186] & 1'b1;
			partial_clause[2][187] 	= partial_clause_prev[2][187] & 1'b1;
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & 1'b1;
			partial_clause[2][190] 	= partial_clause_prev[2][190] & 1'b1;
			partial_clause[2][191] 	= partial_clause_prev[2][191] & 1'b1;
			partial_clause[2][192] 	= partial_clause_prev[2][192] & 1'b1;
			partial_clause[2][193] 	= partial_clause_prev[2][193] & x[19];
			partial_clause[2][194] 	= partial_clause_prev[2][194] & x[44];
			partial_clause[2][195] 	= partial_clause_prev[2][195] & 1'b1;
			partial_clause[2][196] 	= partial_clause_prev[2][196] & 1'b1;
			partial_clause[2][197] 	= partial_clause_prev[2][197] & 1'b1;
			partial_clause[2][198] 	= partial_clause_prev[2][198] & 1'b1;
			partial_clause[2][199] 	= partial_clause_prev[2][199] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & x[42];
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & x[38];
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & x[38];
			partial_clause[3][30] 	= partial_clause_prev[3][30] & x[9];
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & x[36];
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & x[17];
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & x[16];
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[10];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & x[19];
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & x[9];
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & x[40];
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & x[17];
			partial_clause[3][97] 	= partial_clause_prev[3][97] & x[11];
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			partial_clause[3][100] 	= partial_clause_prev[3][100] & ~x[11];
			partial_clause[3][101] 	= partial_clause_prev[3][101] & 1'b1;
			partial_clause[3][102] 	= partial_clause_prev[3][102] & 1'b1;
			partial_clause[3][103] 	= partial_clause_prev[3][103] & 1'b1;
			partial_clause[3][104] 	= partial_clause_prev[3][104] & 1'b1;
			partial_clause[3][105] 	= partial_clause_prev[3][105] & 1'b1;
			partial_clause[3][106] 	= partial_clause_prev[3][106] & ~x[41];
			partial_clause[3][107] 	= partial_clause_prev[3][107] & 1'b1;
			partial_clause[3][108] 	= partial_clause_prev[3][108] & 1'b1;
			partial_clause[3][109] 	= partial_clause_prev[3][109] & 1'b1;
			partial_clause[3][110] 	= partial_clause_prev[3][110] & ~x[40];
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & 1'b1;
			partial_clause[3][113] 	= partial_clause_prev[3][113] & ~x[12] & ~x[39];
			partial_clause[3][114] 	= partial_clause_prev[3][114] & 1'b1;
			partial_clause[3][115] 	= partial_clause_prev[3][115] & 1'b1;
			partial_clause[3][116] 	= partial_clause_prev[3][116] & 1'b1;
			partial_clause[3][117] 	= partial_clause_prev[3][117] & 1'b1;
			partial_clause[3][118] 	= partial_clause_prev[3][118] & 1'b1;
			partial_clause[3][119] 	= partial_clause_prev[3][119] & 1'b1;
			partial_clause[3][120] 	= partial_clause_prev[3][120] & 1'b1;
			partial_clause[3][121] 	= partial_clause_prev[3][121] & 1'b1;
			partial_clause[3][122] 	= partial_clause_prev[3][122] & ~x[42] & ~x[55];
			partial_clause[3][123] 	= partial_clause_prev[3][123] & 1'b1;
			partial_clause[3][124] 	= partial_clause_prev[3][124] & 1'b1;
			partial_clause[3][125] 	= partial_clause_prev[3][125] & 1'b1;
			partial_clause[3][126] 	= partial_clause_prev[3][126] & 1'b1;
			partial_clause[3][127] 	= partial_clause_prev[3][127] & 1'b1;
			partial_clause[3][128] 	= partial_clause_prev[3][128] & 1'b1;
			partial_clause[3][129] 	= partial_clause_prev[3][129] & 1'b1;
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & 1'b1;
			partial_clause[3][132] 	= partial_clause_prev[3][132] & 1'b1;
			partial_clause[3][133] 	= partial_clause_prev[3][133] & 1'b1;
			partial_clause[3][134] 	= partial_clause_prev[3][134] & 1'b1;
			partial_clause[3][135] 	= partial_clause_prev[3][135] & 1'b1;
			partial_clause[3][136] 	= partial_clause_prev[3][136] & 1'b1;
			partial_clause[3][137] 	= partial_clause_prev[3][137] & 1'b1;
			partial_clause[3][138] 	= partial_clause_prev[3][138] & 1'b1;
			partial_clause[3][139] 	= partial_clause_prev[3][139] & 1'b1;
			partial_clause[3][140] 	= partial_clause_prev[3][140] & 1'b1;
			partial_clause[3][141] 	= partial_clause_prev[3][141] & 1'b1;
			partial_clause[3][142] 	= partial_clause_prev[3][142] & 1'b1;
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & 1'b1;
			partial_clause[3][145] 	= partial_clause_prev[3][145] & 1'b1;
			partial_clause[3][146] 	= partial_clause_prev[3][146] & 1'b1;
			partial_clause[3][147] 	= partial_clause_prev[3][147] & 1'b1;
			partial_clause[3][148] 	= partial_clause_prev[3][148] & 1'b1;
			partial_clause[3][149] 	= partial_clause_prev[3][149] & 1'b1;
			partial_clause[3][150] 	= partial_clause_prev[3][150] & 1'b1;
			partial_clause[3][151] 	= partial_clause_prev[3][151] & 1'b1;
			partial_clause[3][152] 	= partial_clause_prev[3][152] & 1'b1;
			partial_clause[3][153] 	= partial_clause_prev[3][153] & 1'b1;
			partial_clause[3][154] 	= partial_clause_prev[3][154] & 1'b1;
			partial_clause[3][155] 	= partial_clause_prev[3][155] & ~x[44];
			partial_clause[3][156] 	= partial_clause_prev[3][156] & ~x[22];
			partial_clause[3][157] 	= partial_clause_prev[3][157] & 1'b1;
			partial_clause[3][158] 	= partial_clause_prev[3][158] & ~x[46];
			partial_clause[3][159] 	= partial_clause_prev[3][159] & 1'b1;
			partial_clause[3][160] 	= partial_clause_prev[3][160] & 1'b1;
			partial_clause[3][161] 	= partial_clause_prev[3][161] & 1'b1;
			partial_clause[3][162] 	= partial_clause_prev[3][162] & 1'b1;
			partial_clause[3][163] 	= partial_clause_prev[3][163] & 1'b1;
			partial_clause[3][164] 	= partial_clause_prev[3][164] & 1'b1;
			partial_clause[3][165] 	= partial_clause_prev[3][165] & 1'b1;
			partial_clause[3][166] 	= partial_clause_prev[3][166] & 1'b1;
			partial_clause[3][167] 	= partial_clause_prev[3][167] & 1'b1;
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & 1'b1;
			partial_clause[3][170] 	= partial_clause_prev[3][170] & 1'b1;
			partial_clause[3][171] 	= partial_clause_prev[3][171] & 1'b1;
			partial_clause[3][172] 	= partial_clause_prev[3][172] & 1'b1;
			partial_clause[3][173] 	= partial_clause_prev[3][173] & 1'b1;
			partial_clause[3][174] 	= partial_clause_prev[3][174] & 1'b1;
			partial_clause[3][175] 	= partial_clause_prev[3][175] & 1'b1;
			partial_clause[3][176] 	= partial_clause_prev[3][176] & 1'b1;
			partial_clause[3][177] 	= partial_clause_prev[3][177] & 1'b1;
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & 1'b1;
			partial_clause[3][180] 	= partial_clause_prev[3][180] & 1'b1;
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & 1'b1;
			partial_clause[3][183] 	= partial_clause_prev[3][183] & ~x[10];
			partial_clause[3][184] 	= partial_clause_prev[3][184] & 1'b1;
			partial_clause[3][185] 	= partial_clause_prev[3][185] & 1'b1;
			partial_clause[3][186] 	= partial_clause_prev[3][186] & 1'b1;
			partial_clause[3][187] 	= partial_clause_prev[3][187] & ~x[42];
			partial_clause[3][188] 	= partial_clause_prev[3][188] & 1'b1;
			partial_clause[3][189] 	= partial_clause_prev[3][189] & 1'b1;
			partial_clause[3][190] 	= partial_clause_prev[3][190] & 1'b1;
			partial_clause[3][191] 	= partial_clause_prev[3][191] & ~x[39];
			partial_clause[3][192] 	= partial_clause_prev[3][192] & 1'b1;
			partial_clause[3][193] 	= partial_clause_prev[3][193] & 1'b1;
			partial_clause[3][194] 	= partial_clause_prev[3][194] & 1'b1;
			partial_clause[3][195] 	= partial_clause_prev[3][195] & 1'b1;
			partial_clause[3][196] 	= partial_clause_prev[3][196] & 1'b1;
			partial_clause[3][197] 	= partial_clause_prev[3][197] & 1'b1;
			partial_clause[3][198] 	= partial_clause_prev[3][198] & 1'b1;
			partial_clause[3][199] 	= partial_clause_prev[3][199] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & x[58];
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & ~x[45];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & x[62];
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & x[58];
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & 1'b1;
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & x[4];
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & 1'b1;
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & x[1];
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & x[31];
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & ~x[15];
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & x[3];
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & x[35];
			partial_clause[4][84] 	= partial_clause_prev[4][84] & x[6];
			partial_clause[4][85] 	= partial_clause_prev[4][85] & ~x[16] & ~x[45];
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			partial_clause[4][100] 	= partial_clause_prev[4][100] & 1'b1;
			partial_clause[4][101] 	= partial_clause_prev[4][101] & 1'b1;
			partial_clause[4][102] 	= partial_clause_prev[4][102] & 1'b1;
			partial_clause[4][103] 	= partial_clause_prev[4][103] & 1'b1;
			partial_clause[4][104] 	= partial_clause_prev[4][104] & 1'b1;
			partial_clause[4][105] 	= partial_clause_prev[4][105] & 1'b1;
			partial_clause[4][106] 	= partial_clause_prev[4][106] & 1'b1;
			partial_clause[4][107] 	= partial_clause_prev[4][107] & 1'b1;
			partial_clause[4][108] 	= partial_clause_prev[4][108] & 1'b1;
			partial_clause[4][109] 	= partial_clause_prev[4][109] & 1'b1;
			partial_clause[4][110] 	= partial_clause_prev[4][110] & 1'b1;
			partial_clause[4][111] 	= partial_clause_prev[4][111] & 1'b1;
			partial_clause[4][112] 	= partial_clause_prev[4][112] & 1'b1;
			partial_clause[4][113] 	= partial_clause_prev[4][113] & 1'b1;
			partial_clause[4][114] 	= partial_clause_prev[4][114] & 1'b1;
			partial_clause[4][115] 	= partial_clause_prev[4][115] & 1'b1;
			partial_clause[4][116] 	= partial_clause_prev[4][116] & 1'b1;
			partial_clause[4][117] 	= partial_clause_prev[4][117] & 1'b1;
			partial_clause[4][118] 	= partial_clause_prev[4][118] & 1'b1;
			partial_clause[4][119] 	= partial_clause_prev[4][119] & 1'b1;
			partial_clause[4][120] 	= partial_clause_prev[4][120] & 1'b1;
			partial_clause[4][121] 	= partial_clause_prev[4][121] & 1'b1;
			partial_clause[4][122] 	= partial_clause_prev[4][122] & 1'b1;
			partial_clause[4][123] 	= partial_clause_prev[4][123] & 1'b1;
			partial_clause[4][124] 	= partial_clause_prev[4][124] & 1'b1;
			partial_clause[4][125] 	= partial_clause_prev[4][125] & 1'b1;
			partial_clause[4][126] 	= partial_clause_prev[4][126] & 1'b1;
			partial_clause[4][127] 	= partial_clause_prev[4][127] & 1'b1;
			partial_clause[4][128] 	= partial_clause_prev[4][128] & 1'b1;
			partial_clause[4][129] 	= partial_clause_prev[4][129] & 1'b1;
			partial_clause[4][130] 	= partial_clause_prev[4][130] & 1'b1;
			partial_clause[4][131] 	= partial_clause_prev[4][131] & 1'b1;
			partial_clause[4][132] 	= partial_clause_prev[4][132] & 1'b1;
			partial_clause[4][133] 	= partial_clause_prev[4][133] & 1'b1;
			partial_clause[4][134] 	= partial_clause_prev[4][134] & 1'b1;
			partial_clause[4][135] 	= partial_clause_prev[4][135] & 1'b1;
			partial_clause[4][136] 	= partial_clause_prev[4][136] & 1'b1;
			partial_clause[4][137] 	= partial_clause_prev[4][137] & 1'b1;
			partial_clause[4][138] 	= partial_clause_prev[4][138] & 1'b1;
			partial_clause[4][139] 	= partial_clause_prev[4][139] & 1'b1;
			partial_clause[4][140] 	= partial_clause_prev[4][140] & 1'b1;
			partial_clause[4][141] 	= partial_clause_prev[4][141] & 1'b1;
			partial_clause[4][142] 	= partial_clause_prev[4][142] & 1'b1;
			partial_clause[4][143] 	= partial_clause_prev[4][143] & 1'b1;
			partial_clause[4][144] 	= partial_clause_prev[4][144] & 1'b1;
			partial_clause[4][145] 	= partial_clause_prev[4][145] & 1'b1;
			partial_clause[4][146] 	= partial_clause_prev[4][146] & 1'b1;
			partial_clause[4][147] 	= partial_clause_prev[4][147] & 1'b1;
			partial_clause[4][148] 	= partial_clause_prev[4][148] & 1'b1;
			partial_clause[4][149] 	= partial_clause_prev[4][149] & 1'b1;
			partial_clause[4][150] 	= partial_clause_prev[4][150] & 1'b1;
			partial_clause[4][151] 	= partial_clause_prev[4][151] & 1'b1;
			partial_clause[4][152] 	= partial_clause_prev[4][152] & 1'b1;
			partial_clause[4][153] 	= partial_clause_prev[4][153] & 1'b1;
			partial_clause[4][154] 	= partial_clause_prev[4][154] & 1'b1;
			partial_clause[4][155] 	= partial_clause_prev[4][155] & 1'b1;
			partial_clause[4][156] 	= partial_clause_prev[4][156] & 1'b1;
			partial_clause[4][157] 	= partial_clause_prev[4][157] & ~x[58];
			partial_clause[4][158] 	= partial_clause_prev[4][158] & 1'b1;
			partial_clause[4][159] 	= partial_clause_prev[4][159] & 1'b1;
			partial_clause[4][160] 	= partial_clause_prev[4][160] & 1'b1;
			partial_clause[4][161] 	= partial_clause_prev[4][161] & ~x[33] & ~x[60];
			partial_clause[4][162] 	= partial_clause_prev[4][162] & 1'b1;
			partial_clause[4][163] 	= partial_clause_prev[4][163] & ~x[14];
			partial_clause[4][164] 	= partial_clause_prev[4][164] & 1'b1;
			partial_clause[4][165] 	= partial_clause_prev[4][165] & 1'b1;
			partial_clause[4][166] 	= partial_clause_prev[4][166] & 1'b1;
			partial_clause[4][167] 	= partial_clause_prev[4][167] & 1'b1;
			partial_clause[4][168] 	= partial_clause_prev[4][168] & 1'b1;
			partial_clause[4][169] 	= partial_clause_prev[4][169] & 1'b1;
			partial_clause[4][170] 	= partial_clause_prev[4][170] & 1'b1;
			partial_clause[4][171] 	= partial_clause_prev[4][171] & 1'b1;
			partial_clause[4][172] 	= partial_clause_prev[4][172] & 1'b1;
			partial_clause[4][173] 	= partial_clause_prev[4][173] & 1'b1;
			partial_clause[4][174] 	= partial_clause_prev[4][174] & 1'b1;
			partial_clause[4][175] 	= partial_clause_prev[4][175] & 1'b1;
			partial_clause[4][176] 	= partial_clause_prev[4][176] & 1'b1;
			partial_clause[4][177] 	= partial_clause_prev[4][177] & 1'b1;
			partial_clause[4][178] 	= partial_clause_prev[4][178] & 1'b1;
			partial_clause[4][179] 	= partial_clause_prev[4][179] & 1'b1;
			partial_clause[4][180] 	= partial_clause_prev[4][180] & 1'b1;
			partial_clause[4][181] 	= partial_clause_prev[4][181] & 1'b1;
			partial_clause[4][182] 	= partial_clause_prev[4][182] & 1'b1;
			partial_clause[4][183] 	= partial_clause_prev[4][183] & 1'b1;
			partial_clause[4][184] 	= partial_clause_prev[4][184] & 1'b1;
			partial_clause[4][185] 	= partial_clause_prev[4][185] & 1'b1;
			partial_clause[4][186] 	= partial_clause_prev[4][186] & 1'b1;
			partial_clause[4][187] 	= partial_clause_prev[4][187] & 1'b1;
			partial_clause[4][188] 	= partial_clause_prev[4][188] & ~x[12];
			partial_clause[4][189] 	= partial_clause_prev[4][189] & ~x[51];
			partial_clause[4][190] 	= partial_clause_prev[4][190] & 1'b1;
			partial_clause[4][191] 	= partial_clause_prev[4][191] & 1'b1;
			partial_clause[4][192] 	= partial_clause_prev[4][192] & 1'b1;
			partial_clause[4][193] 	= partial_clause_prev[4][193] & 1'b1;
			partial_clause[4][194] 	= partial_clause_prev[4][194] & 1'b1;
			partial_clause[4][195] 	= partial_clause_prev[4][195] & 1'b1;
			partial_clause[4][196] 	= partial_clause_prev[4][196] & 1'b1;
			partial_clause[4][197] 	= partial_clause_prev[4][197] & 1'b1;
			partial_clause[4][198] 	= partial_clause_prev[4][198] & 1'b1;
			partial_clause[4][199] 	= partial_clause_prev[4][199] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & x[15];
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & x[54];
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & x[17];
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & x[53];
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & ~x[11];
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & x[18];
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & x[19];
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			partial_clause[5][100] 	= partial_clause_prev[5][100] & 1'b1;
			partial_clause[5][101] 	= partial_clause_prev[5][101] & 1'b1;
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & 1'b1;
			partial_clause[5][104] 	= partial_clause_prev[5][104] & 1'b1;
			partial_clause[5][105] 	= partial_clause_prev[5][105] & 1'b1;
			partial_clause[5][106] 	= partial_clause_prev[5][106] & 1'b1;
			partial_clause[5][107] 	= partial_clause_prev[5][107] & 1'b1;
			partial_clause[5][108] 	= partial_clause_prev[5][108] & 1'b1;
			partial_clause[5][109] 	= partial_clause_prev[5][109] & 1'b1;
			partial_clause[5][110] 	= partial_clause_prev[5][110] & 1'b1;
			partial_clause[5][111] 	= partial_clause_prev[5][111] & 1'b1;
			partial_clause[5][112] 	= partial_clause_prev[5][112] & 1'b1;
			partial_clause[5][113] 	= partial_clause_prev[5][113] & 1'b1;
			partial_clause[5][114] 	= partial_clause_prev[5][114] & 1'b1;
			partial_clause[5][115] 	= partial_clause_prev[5][115] & 1'b1;
			partial_clause[5][116] 	= partial_clause_prev[5][116] & 1'b1;
			partial_clause[5][117] 	= partial_clause_prev[5][117] & 1'b1;
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & 1'b1;
			partial_clause[5][120] 	= partial_clause_prev[5][120] & 1'b1;
			partial_clause[5][121] 	= partial_clause_prev[5][121] & 1'b1;
			partial_clause[5][122] 	= partial_clause_prev[5][122] & 1'b1;
			partial_clause[5][123] 	= partial_clause_prev[5][123] & 1'b1;
			partial_clause[5][124] 	= partial_clause_prev[5][124] & 1'b1;
			partial_clause[5][125] 	= partial_clause_prev[5][125] & 1'b1;
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & 1'b1;
			partial_clause[5][128] 	= partial_clause_prev[5][128] & 1'b1;
			partial_clause[5][129] 	= partial_clause_prev[5][129] & 1'b1;
			partial_clause[5][130] 	= partial_clause_prev[5][130] & ~x[21];
			partial_clause[5][131] 	= partial_clause_prev[5][131] & 1'b1;
			partial_clause[5][132] 	= partial_clause_prev[5][132] & 1'b1;
			partial_clause[5][133] 	= partial_clause_prev[5][133] & 1'b1;
			partial_clause[5][134] 	= partial_clause_prev[5][134] & 1'b1;
			partial_clause[5][135] 	= partial_clause_prev[5][135] & 1'b1;
			partial_clause[5][136] 	= partial_clause_prev[5][136] & 1'b1;
			partial_clause[5][137] 	= partial_clause_prev[5][137] & 1'b1;
			partial_clause[5][138] 	= partial_clause_prev[5][138] & 1'b1;
			partial_clause[5][139] 	= partial_clause_prev[5][139] & 1'b1;
			partial_clause[5][140] 	= partial_clause_prev[5][140] & 1'b1;
			partial_clause[5][141] 	= partial_clause_prev[5][141] & 1'b1;
			partial_clause[5][142] 	= partial_clause_prev[5][142] & 1'b1;
			partial_clause[5][143] 	= partial_clause_prev[5][143] & 1'b1;
			partial_clause[5][144] 	= partial_clause_prev[5][144] & 1'b1;
			partial_clause[5][145] 	= partial_clause_prev[5][145] & 1'b1;
			partial_clause[5][146] 	= partial_clause_prev[5][146] & 1'b1;
			partial_clause[5][147] 	= partial_clause_prev[5][147] & 1'b1;
			partial_clause[5][148] 	= partial_clause_prev[5][148] & 1'b1;
			partial_clause[5][149] 	= partial_clause_prev[5][149] & 1'b1;
			partial_clause[5][150] 	= partial_clause_prev[5][150] & 1'b1;
			partial_clause[5][151] 	= partial_clause_prev[5][151] & 1'b1;
			partial_clause[5][152] 	= partial_clause_prev[5][152] & 1'b1;
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & 1'b1;
			partial_clause[5][155] 	= partial_clause_prev[5][155] & x[4];
			partial_clause[5][156] 	= partial_clause_prev[5][156] & 1'b1;
			partial_clause[5][157] 	= partial_clause_prev[5][157] & 1'b1;
			partial_clause[5][158] 	= partial_clause_prev[5][158] & 1'b1;
			partial_clause[5][159] 	= partial_clause_prev[5][159] & 1'b1;
			partial_clause[5][160] 	= partial_clause_prev[5][160] & 1'b1;
			partial_clause[5][161] 	= partial_clause_prev[5][161] & 1'b1;
			partial_clause[5][162] 	= partial_clause_prev[5][162] & 1'b1;
			partial_clause[5][163] 	= partial_clause_prev[5][163] & 1'b1;
			partial_clause[5][164] 	= partial_clause_prev[5][164] & 1'b1;
			partial_clause[5][165] 	= partial_clause_prev[5][165] & 1'b1;
			partial_clause[5][166] 	= partial_clause_prev[5][166] & 1'b1;
			partial_clause[5][167] 	= partial_clause_prev[5][167] & 1'b1;
			partial_clause[5][168] 	= partial_clause_prev[5][168] & 1'b1;
			partial_clause[5][169] 	= partial_clause_prev[5][169] & 1'b1;
			partial_clause[5][170] 	= partial_clause_prev[5][170] & 1'b1;
			partial_clause[5][171] 	= partial_clause_prev[5][171] & 1'b1;
			partial_clause[5][172] 	= partial_clause_prev[5][172] & 1'b1;
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & 1'b1;
			partial_clause[5][175] 	= partial_clause_prev[5][175] & 1'b1;
			partial_clause[5][176] 	= partial_clause_prev[5][176] & 1'b1;
			partial_clause[5][177] 	= partial_clause_prev[5][177] & 1'b1;
			partial_clause[5][178] 	= partial_clause_prev[5][178] & 1'b1;
			partial_clause[5][179] 	= partial_clause_prev[5][179] & 1'b1;
			partial_clause[5][180] 	= partial_clause_prev[5][180] & 1'b1;
			partial_clause[5][181] 	= partial_clause_prev[5][181] & 1'b1;
			partial_clause[5][182] 	= partial_clause_prev[5][182] & 1'b1;
			partial_clause[5][183] 	= partial_clause_prev[5][183] & 1'b1;
			partial_clause[5][184] 	= partial_clause_prev[5][184] & 1'b1;
			partial_clause[5][185] 	= partial_clause_prev[5][185] & 1'b1;
			partial_clause[5][186] 	= partial_clause_prev[5][186] & 1'b1;
			partial_clause[5][187] 	= partial_clause_prev[5][187] & 1'b1;
			partial_clause[5][188] 	= partial_clause_prev[5][188] & 1'b1;
			partial_clause[5][189] 	= partial_clause_prev[5][189] & 1'b1;
			partial_clause[5][190] 	= partial_clause_prev[5][190] & 1'b1;
			partial_clause[5][191] 	= partial_clause_prev[5][191] & 1'b1;
			partial_clause[5][192] 	= partial_clause_prev[5][192] & 1'b1;
			partial_clause[5][193] 	= partial_clause_prev[5][193] & 1'b1;
			partial_clause[5][194] 	= partial_clause_prev[5][194] & 1'b1;
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & 1'b1;
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & 1'b1;
			partial_clause[5][199] 	= partial_clause_prev[5][199] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & ~x[47];
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & ~x[19];
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & ~x[16];
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & ~x[16];
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & ~x[21];
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & ~x[18];
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & ~x[14] & ~x[18];
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			partial_clause[6][100] 	= partial_clause_prev[6][100] & 1'b1;
			partial_clause[6][101] 	= partial_clause_prev[6][101] & 1'b1;
			partial_clause[6][102] 	= partial_clause_prev[6][102] & 1'b1;
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & x[17];
			partial_clause[6][105] 	= partial_clause_prev[6][105] & 1'b1;
			partial_clause[6][106] 	= partial_clause_prev[6][106] & 1'b1;
			partial_clause[6][107] 	= partial_clause_prev[6][107] & 1'b1;
			partial_clause[6][108] 	= partial_clause_prev[6][108] & 1'b1;
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & 1'b1;
			partial_clause[6][111] 	= partial_clause_prev[6][111] & 1'b1;
			partial_clause[6][112] 	= partial_clause_prev[6][112] & 1'b1;
			partial_clause[6][113] 	= partial_clause_prev[6][113] & 1'b1;
			partial_clause[6][114] 	= partial_clause_prev[6][114] & x[12];
			partial_clause[6][115] 	= partial_clause_prev[6][115] & 1'b1;
			partial_clause[6][116] 	= partial_clause_prev[6][116] & 1'b1;
			partial_clause[6][117] 	= partial_clause_prev[6][117] & 1'b1;
			partial_clause[6][118] 	= partial_clause_prev[6][118] & 1'b1;
			partial_clause[6][119] 	= partial_clause_prev[6][119] & 1'b1;
			partial_clause[6][120] 	= partial_clause_prev[6][120] & 1'b1;
			partial_clause[6][121] 	= partial_clause_prev[6][121] & 1'b1;
			partial_clause[6][122] 	= partial_clause_prev[6][122] & 1'b1;
			partial_clause[6][123] 	= partial_clause_prev[6][123] & 1'b1;
			partial_clause[6][124] 	= partial_clause_prev[6][124] & x[44];
			partial_clause[6][125] 	= partial_clause_prev[6][125] & 1'b1;
			partial_clause[6][126] 	= partial_clause_prev[6][126] & 1'b1;
			partial_clause[6][127] 	= partial_clause_prev[6][127] & x[44];
			partial_clause[6][128] 	= partial_clause_prev[6][128] & x[48];
			partial_clause[6][129] 	= partial_clause_prev[6][129] & 1'b1;
			partial_clause[6][130] 	= partial_clause_prev[6][130] & 1'b1;
			partial_clause[6][131] 	= partial_clause_prev[6][131] & 1'b1;
			partial_clause[6][132] 	= partial_clause_prev[6][132] & 1'b1;
			partial_clause[6][133] 	= partial_clause_prev[6][133] & 1'b1;
			partial_clause[6][134] 	= partial_clause_prev[6][134] & 1'b1;
			partial_clause[6][135] 	= partial_clause_prev[6][135] & 1'b1;
			partial_clause[6][136] 	= partial_clause_prev[6][136] & ~x[48];
			partial_clause[6][137] 	= partial_clause_prev[6][137] & 1'b1;
			partial_clause[6][138] 	= partial_clause_prev[6][138] & 1'b1;
			partial_clause[6][139] 	= partial_clause_prev[6][139] & 1'b1;
			partial_clause[6][140] 	= partial_clause_prev[6][140] & 1'b1;
			partial_clause[6][141] 	= partial_clause_prev[6][141] & 1'b1;
			partial_clause[6][142] 	= partial_clause_prev[6][142] & 1'b1;
			partial_clause[6][143] 	= partial_clause_prev[6][143] & 1'b1;
			partial_clause[6][144] 	= partial_clause_prev[6][144] & 1'b1;
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & ~x[23];
			partial_clause[6][147] 	= partial_clause_prev[6][147] & 1'b1;
			partial_clause[6][148] 	= partial_clause_prev[6][148] & x[46];
			partial_clause[6][149] 	= partial_clause_prev[6][149] & 1'b1;
			partial_clause[6][150] 	= partial_clause_prev[6][150] & 1'b1;
			partial_clause[6][151] 	= partial_clause_prev[6][151] & 1'b1;
			partial_clause[6][152] 	= partial_clause_prev[6][152] & 1'b1;
			partial_clause[6][153] 	= partial_clause_prev[6][153] & 1'b1;
			partial_clause[6][154] 	= partial_clause_prev[6][154] & 1'b1;
			partial_clause[6][155] 	= partial_clause_prev[6][155] & 1'b1;
			partial_clause[6][156] 	= partial_clause_prev[6][156] & 1'b1;
			partial_clause[6][157] 	= partial_clause_prev[6][157] & 1'b1;
			partial_clause[6][158] 	= partial_clause_prev[6][158] & 1'b1;
			partial_clause[6][159] 	= partial_clause_prev[6][159] & x[20];
			partial_clause[6][160] 	= partial_clause_prev[6][160] & 1'b1;
			partial_clause[6][161] 	= partial_clause_prev[6][161] & x[13];
			partial_clause[6][162] 	= partial_clause_prev[6][162] & 1'b1;
			partial_clause[6][163] 	= partial_clause_prev[6][163] & 1'b1;
			partial_clause[6][164] 	= partial_clause_prev[6][164] & x[41];
			partial_clause[6][165] 	= partial_clause_prev[6][165] & 1'b1;
			partial_clause[6][166] 	= partial_clause_prev[6][166] & 1'b1;
			partial_clause[6][167] 	= partial_clause_prev[6][167] & 1'b1;
			partial_clause[6][168] 	= partial_clause_prev[6][168] & 1'b1;
			partial_clause[6][169] 	= partial_clause_prev[6][169] & 1'b1;
			partial_clause[6][170] 	= partial_clause_prev[6][170] & 1'b1;
			partial_clause[6][171] 	= partial_clause_prev[6][171] & 1'b1;
			partial_clause[6][172] 	= partial_clause_prev[6][172] & 1'b1;
			partial_clause[6][173] 	= partial_clause_prev[6][173] & 1'b1;
			partial_clause[6][174] 	= partial_clause_prev[6][174] & 1'b1;
			partial_clause[6][175] 	= partial_clause_prev[6][175] & 1'b1;
			partial_clause[6][176] 	= partial_clause_prev[6][176] & 1'b1;
			partial_clause[6][177] 	= partial_clause_prev[6][177] & 1'b1;
			partial_clause[6][178] 	= partial_clause_prev[6][178] & 1'b1;
			partial_clause[6][179] 	= partial_clause_prev[6][179] & 1'b1;
			partial_clause[6][180] 	= partial_clause_prev[6][180] & 1'b1;
			partial_clause[6][181] 	= partial_clause_prev[6][181] & 1'b1;
			partial_clause[6][182] 	= partial_clause_prev[6][182] & 1'b1;
			partial_clause[6][183] 	= partial_clause_prev[6][183] & 1'b1;
			partial_clause[6][184] 	= partial_clause_prev[6][184] & 1'b1;
			partial_clause[6][185] 	= partial_clause_prev[6][185] & 1'b1;
			partial_clause[6][186] 	= partial_clause_prev[6][186] & 1'b1;
			partial_clause[6][187] 	= partial_clause_prev[6][187] & 1'b1;
			partial_clause[6][188] 	= partial_clause_prev[6][188] & x[14];
			partial_clause[6][189] 	= partial_clause_prev[6][189] & 1'b1;
			partial_clause[6][190] 	= partial_clause_prev[6][190] & 1'b1;
			partial_clause[6][191] 	= partial_clause_prev[6][191] & 1'b1;
			partial_clause[6][192] 	= partial_clause_prev[6][192] & x[15];
			partial_clause[6][193] 	= partial_clause_prev[6][193] & 1'b1;
			partial_clause[6][194] 	= partial_clause_prev[6][194] & 1'b1;
			partial_clause[6][195] 	= partial_clause_prev[6][195] & x[46];
			partial_clause[6][196] 	= partial_clause_prev[6][196] & 1'b1;
			partial_clause[6][197] 	= partial_clause_prev[6][197] & 1'b1;
			partial_clause[6][198] 	= partial_clause_prev[6][198] & 1'b1;
			partial_clause[6][199] 	= partial_clause_prev[6][199] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & ~x[22];
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & x[29];
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & x[37];
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & x[38];
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & x[58];
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & ~x[19] & x[42];
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & x[36];
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & x[40];
			partial_clause[7][74] 	= partial_clause_prev[7][74] & x[38];
			partial_clause[7][75] 	= partial_clause_prev[7][75] & ~x[15] & ~x[42] & ~x[43] & x[46];
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & x[45];
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & ~x[51];
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			partial_clause[7][100] 	= partial_clause_prev[7][100] & 1'b1;
			partial_clause[7][101] 	= partial_clause_prev[7][101] & 1'b1;
			partial_clause[7][102] 	= partial_clause_prev[7][102] & 1'b1;
			partial_clause[7][103] 	= partial_clause_prev[7][103] & 1'b1;
			partial_clause[7][104] 	= partial_clause_prev[7][104] & 1'b1;
			partial_clause[7][105] 	= partial_clause_prev[7][105] & 1'b1;
			partial_clause[7][106] 	= partial_clause_prev[7][106] & 1'b1;
			partial_clause[7][107] 	= partial_clause_prev[7][107] & 1'b1;
			partial_clause[7][108] 	= partial_clause_prev[7][108] & ~x[39];
			partial_clause[7][109] 	= partial_clause_prev[7][109] & 1'b1;
			partial_clause[7][110] 	= partial_clause_prev[7][110] & 1'b1;
			partial_clause[7][111] 	= partial_clause_prev[7][111] & 1'b1;
			partial_clause[7][112] 	= partial_clause_prev[7][112] & 1'b1;
			partial_clause[7][113] 	= partial_clause_prev[7][113] & 1'b1;
			partial_clause[7][114] 	= partial_clause_prev[7][114] & 1'b1;
			partial_clause[7][115] 	= partial_clause_prev[7][115] & 1'b1;
			partial_clause[7][116] 	= partial_clause_prev[7][116] & 1'b1;
			partial_clause[7][117] 	= partial_clause_prev[7][117] & 1'b1;
			partial_clause[7][118] 	= partial_clause_prev[7][118] & 1'b1;
			partial_clause[7][119] 	= partial_clause_prev[7][119] & 1'b1;
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & 1'b1;
			partial_clause[7][123] 	= partial_clause_prev[7][123] & 1'b1;
			partial_clause[7][124] 	= partial_clause_prev[7][124] & 1'b1;
			partial_clause[7][125] 	= partial_clause_prev[7][125] & 1'b1;
			partial_clause[7][126] 	= partial_clause_prev[7][126] & 1'b1;
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & 1'b1;
			partial_clause[7][129] 	= partial_clause_prev[7][129] & 1'b1;
			partial_clause[7][130] 	= partial_clause_prev[7][130] & 1'b1;
			partial_clause[7][131] 	= partial_clause_prev[7][131] & 1'b1;
			partial_clause[7][132] 	= partial_clause_prev[7][132] & 1'b1;
			partial_clause[7][133] 	= partial_clause_prev[7][133] & 1'b1;
			partial_clause[7][134] 	= partial_clause_prev[7][134] & 1'b1;
			partial_clause[7][135] 	= partial_clause_prev[7][135] & 1'b1;
			partial_clause[7][136] 	= partial_clause_prev[7][136] & 1'b1;
			partial_clause[7][137] 	= partial_clause_prev[7][137] & 1'b1;
			partial_clause[7][138] 	= partial_clause_prev[7][138] & 1'b1;
			partial_clause[7][139] 	= partial_clause_prev[7][139] & 1'b1;
			partial_clause[7][140] 	= partial_clause_prev[7][140] & 1'b1;
			partial_clause[7][141] 	= partial_clause_prev[7][141] & 1'b1;
			partial_clause[7][142] 	= partial_clause_prev[7][142] & 1'b1;
			partial_clause[7][143] 	= partial_clause_prev[7][143] & 1'b1;
			partial_clause[7][144] 	= partial_clause_prev[7][144] & 1'b1;
			partial_clause[7][145] 	= partial_clause_prev[7][145] & 1'b1;
			partial_clause[7][146] 	= partial_clause_prev[7][146] & 1'b1;
			partial_clause[7][147] 	= partial_clause_prev[7][147] & 1'b1;
			partial_clause[7][148] 	= partial_clause_prev[7][148] & 1'b1;
			partial_clause[7][149] 	= partial_clause_prev[7][149] & 1'b1;
			partial_clause[7][150] 	= partial_clause_prev[7][150] & 1'b1;
			partial_clause[7][151] 	= partial_clause_prev[7][151] & 1'b1;
			partial_clause[7][152] 	= partial_clause_prev[7][152] & 1'b1;
			partial_clause[7][153] 	= partial_clause_prev[7][153] & 1'b1;
			partial_clause[7][154] 	= partial_clause_prev[7][154] & 1'b1;
			partial_clause[7][155] 	= partial_clause_prev[7][155] & 1'b1;
			partial_clause[7][156] 	= partial_clause_prev[7][156] & 1'b1;
			partial_clause[7][157] 	= partial_clause_prev[7][157] & 1'b1;
			partial_clause[7][158] 	= partial_clause_prev[7][158] & 1'b1;
			partial_clause[7][159] 	= partial_clause_prev[7][159] & 1'b1;
			partial_clause[7][160] 	= partial_clause_prev[7][160] & 1'b1;
			partial_clause[7][161] 	= partial_clause_prev[7][161] & 1'b1;
			partial_clause[7][162] 	= partial_clause_prev[7][162] & 1'b1;
			partial_clause[7][163] 	= partial_clause_prev[7][163] & 1'b1;
			partial_clause[7][164] 	= partial_clause_prev[7][164] & 1'b1;
			partial_clause[7][165] 	= partial_clause_prev[7][165] & 1'b1;
			partial_clause[7][166] 	= partial_clause_prev[7][166] & 1'b1;
			partial_clause[7][167] 	= partial_clause_prev[7][167] & 1'b1;
			partial_clause[7][168] 	= partial_clause_prev[7][168] & 1'b1;
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & 1'b1;
			partial_clause[7][171] 	= partial_clause_prev[7][171] & ~x[1];
			partial_clause[7][172] 	= partial_clause_prev[7][172] & 1'b1;
			partial_clause[7][173] 	= partial_clause_prev[7][173] & 1'b1;
			partial_clause[7][174] 	= partial_clause_prev[7][174] & 1'b1;
			partial_clause[7][175] 	= partial_clause_prev[7][175] & ~x[38];
			partial_clause[7][176] 	= partial_clause_prev[7][176] & 1'b1;
			partial_clause[7][177] 	= partial_clause_prev[7][177] & 1'b1;
			partial_clause[7][178] 	= partial_clause_prev[7][178] & 1'b1;
			partial_clause[7][179] 	= partial_clause_prev[7][179] & 1'b1;
			partial_clause[7][180] 	= partial_clause_prev[7][180] & 1'b1;
			partial_clause[7][181] 	= partial_clause_prev[7][181] & 1'b1;
			partial_clause[7][182] 	= partial_clause_prev[7][182] & 1'b1;
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & 1'b1;
			partial_clause[7][185] 	= partial_clause_prev[7][185] & 1'b1;
			partial_clause[7][186] 	= partial_clause_prev[7][186] & ~x[37];
			partial_clause[7][187] 	= partial_clause_prev[7][187] & 1'b1;
			partial_clause[7][188] 	= partial_clause_prev[7][188] & 1'b1;
			partial_clause[7][189] 	= partial_clause_prev[7][189] & 1'b1;
			partial_clause[7][190] 	= partial_clause_prev[7][190] & 1'b1;
			partial_clause[7][191] 	= partial_clause_prev[7][191] & 1'b1;
			partial_clause[7][192] 	= partial_clause_prev[7][192] & 1'b1;
			partial_clause[7][193] 	= partial_clause_prev[7][193] & 1'b1;
			partial_clause[7][194] 	= partial_clause_prev[7][194] & 1'b1;
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & ~x[32];
			partial_clause[7][197] 	= partial_clause_prev[7][197] & 1'b1;
			partial_clause[7][198] 	= partial_clause_prev[7][198] & 1'b1;
			partial_clause[7][199] 	= partial_clause_prev[7][199] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & x[22];
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & x[20];
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & x[47];
			partial_clause[8][10] 	= partial_clause_prev[8][10] & x[16];
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & x[16];
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & ~x[11] & x[18];
			partial_clause[8][25] 	= partial_clause_prev[8][25] & x[19];
			partial_clause[8][26] 	= partial_clause_prev[8][26] & x[17];
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & x[17];
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & x[0];
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & x[15];
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & x[19];
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & x[20];
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & x[6];
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & x[31];
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & x[17];
			partial_clause[8][57] 	= partial_clause_prev[8][57] & x[19];
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & x[17];
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & x[51];
			partial_clause[8][75] 	= partial_clause_prev[8][75] & x[61];
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & x[18];
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & x[18];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & x[15];
			partial_clause[8][92] 	= partial_clause_prev[8][92] & x[23];
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & x[15];
			partial_clause[8][95] 	= partial_clause_prev[8][95] & x[13];
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			partial_clause[8][100] 	= partial_clause_prev[8][100] & 1'b1;
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & 1'b1;
			partial_clause[8][103] 	= partial_clause_prev[8][103] & 1'b1;
			partial_clause[8][104] 	= partial_clause_prev[8][104] & 1'b1;
			partial_clause[8][105] 	= partial_clause_prev[8][105] & 1'b1;
			partial_clause[8][106] 	= partial_clause_prev[8][106] & 1'b1;
			partial_clause[8][107] 	= partial_clause_prev[8][107] & 1'b1;
			partial_clause[8][108] 	= partial_clause_prev[8][108] & 1'b1;
			partial_clause[8][109] 	= partial_clause_prev[8][109] & 1'b1;
			partial_clause[8][110] 	= partial_clause_prev[8][110] & 1'b1;
			partial_clause[8][111] 	= partial_clause_prev[8][111] & 1'b1;
			partial_clause[8][112] 	= partial_clause_prev[8][112] & 1'b1;
			partial_clause[8][113] 	= partial_clause_prev[8][113] & 1'b1;
			partial_clause[8][114] 	= partial_clause_prev[8][114] & 1'b1;
			partial_clause[8][115] 	= partial_clause_prev[8][115] & 1'b1;
			partial_clause[8][116] 	= partial_clause_prev[8][116] & 1'b1;
			partial_clause[8][117] 	= partial_clause_prev[8][117] & 1'b1;
			partial_clause[8][118] 	= partial_clause_prev[8][118] & 1'b1;
			partial_clause[8][119] 	= partial_clause_prev[8][119] & 1'b1;
			partial_clause[8][120] 	= partial_clause_prev[8][120] & 1'b1;
			partial_clause[8][121] 	= partial_clause_prev[8][121] & 1'b1;
			partial_clause[8][122] 	= partial_clause_prev[8][122] & 1'b1;
			partial_clause[8][123] 	= partial_clause_prev[8][123] & 1'b1;
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & x[28];
			partial_clause[8][126] 	= partial_clause_prev[8][126] & 1'b1;
			partial_clause[8][127] 	= partial_clause_prev[8][127] & ~x[21] & ~x[23];
			partial_clause[8][128] 	= partial_clause_prev[8][128] & 1'b1;
			partial_clause[8][129] 	= partial_clause_prev[8][129] & 1'b1;
			partial_clause[8][130] 	= partial_clause_prev[8][130] & 1'b1;
			partial_clause[8][131] 	= partial_clause_prev[8][131] & 1'b1;
			partial_clause[8][132] 	= partial_clause_prev[8][132] & 1'b1;
			partial_clause[8][133] 	= partial_clause_prev[8][133] & 1'b1;
			partial_clause[8][134] 	= partial_clause_prev[8][134] & 1'b1;
			partial_clause[8][135] 	= partial_clause_prev[8][135] & ~x[44] & ~x[45];
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & 1'b1;
			partial_clause[8][138] 	= partial_clause_prev[8][138] & x[29];
			partial_clause[8][139] 	= partial_clause_prev[8][139] & 1'b1;
			partial_clause[8][140] 	= partial_clause_prev[8][140] & 1'b1;
			partial_clause[8][141] 	= partial_clause_prev[8][141] & ~x[15] & ~x[16];
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & 1'b1;
			partial_clause[8][144] 	= partial_clause_prev[8][144] & 1'b1;
			partial_clause[8][145] 	= partial_clause_prev[8][145] & 1'b1;
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & 1'b1;
			partial_clause[8][148] 	= partial_clause_prev[8][148] & 1'b1;
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & 1'b1;
			partial_clause[8][151] 	= partial_clause_prev[8][151] & 1'b1;
			partial_clause[8][152] 	= partial_clause_prev[8][152] & 1'b1;
			partial_clause[8][153] 	= partial_clause_prev[8][153] & 1'b1;
			partial_clause[8][154] 	= partial_clause_prev[8][154] & 1'b1;
			partial_clause[8][155] 	= partial_clause_prev[8][155] & 1'b1;
			partial_clause[8][156] 	= partial_clause_prev[8][156] & 1'b1;
			partial_clause[8][157] 	= partial_clause_prev[8][157] & 1'b1;
			partial_clause[8][158] 	= partial_clause_prev[8][158] & 1'b1;
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & 1'b1;
			partial_clause[8][161] 	= partial_clause_prev[8][161] & x[63];
			partial_clause[8][162] 	= partial_clause_prev[8][162] & 1'b1;
			partial_clause[8][163] 	= partial_clause_prev[8][163] & ~x[47];
			partial_clause[8][164] 	= partial_clause_prev[8][164] & 1'b1;
			partial_clause[8][165] 	= partial_clause_prev[8][165] & ~x[15] & ~x[23] & ~x[41];
			partial_clause[8][166] 	= partial_clause_prev[8][166] & 1'b1;
			partial_clause[8][167] 	= partial_clause_prev[8][167] & 1'b1;
			partial_clause[8][168] 	= partial_clause_prev[8][168] & 1'b1;
			partial_clause[8][169] 	= partial_clause_prev[8][169] & 1'b1;
			partial_clause[8][170] 	= partial_clause_prev[8][170] & 1'b1;
			partial_clause[8][171] 	= partial_clause_prev[8][171] & 1'b1;
			partial_clause[8][172] 	= partial_clause_prev[8][172] & 1'b1;
			partial_clause[8][173] 	= partial_clause_prev[8][173] & 1'b1;
			partial_clause[8][174] 	= partial_clause_prev[8][174] & 1'b1;
			partial_clause[8][175] 	= partial_clause_prev[8][175] & 1'b1;
			partial_clause[8][176] 	= partial_clause_prev[8][176] & 1'b1;
			partial_clause[8][177] 	= partial_clause_prev[8][177] & 1'b1;
			partial_clause[8][178] 	= partial_clause_prev[8][178] & 1'b1;
			partial_clause[8][179] 	= partial_clause_prev[8][179] & ~x[12] & ~x[21] & ~x[47];
			partial_clause[8][180] 	= partial_clause_prev[8][180] & 1'b1;
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & 1'b1;
			partial_clause[8][183] 	= partial_clause_prev[8][183] & 1'b1;
			partial_clause[8][184] 	= partial_clause_prev[8][184] & 1'b1;
			partial_clause[8][185] 	= partial_clause_prev[8][185] & x[55];
			partial_clause[8][186] 	= partial_clause_prev[8][186] & 1'b1;
			partial_clause[8][187] 	= partial_clause_prev[8][187] & 1'b1;
			partial_clause[8][188] 	= partial_clause_prev[8][188] & 1'b1;
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & ~x[48];
			partial_clause[8][191] 	= partial_clause_prev[8][191] & 1'b1;
			partial_clause[8][192] 	= partial_clause_prev[8][192] & 1'b1;
			partial_clause[8][193] 	= partial_clause_prev[8][193] & 1'b1;
			partial_clause[8][194] 	= partial_clause_prev[8][194] & ~x[12];
			partial_clause[8][195] 	= partial_clause_prev[8][195] & ~x[20];
			partial_clause[8][196] 	= partial_clause_prev[8][196] & 1'b1;
			partial_clause[8][197] 	= partial_clause_prev[8][197] & 1'b1;
			partial_clause[8][198] 	= partial_clause_prev[8][198] & 1'b1;
			partial_clause[8][199] 	= partial_clause_prev[8][199] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & x[58];
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & ~x[60];
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & x[57];
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & x[55];
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & x[53];
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & x[26];
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & ~x[15];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & ~x[42];
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & x[52];
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & x[27];
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & x[27];
			partial_clause[9][51] 	= partial_clause_prev[9][51] & x[62];
			partial_clause[9][52] 	= partial_clause_prev[9][52] & x[32];
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & x[57];
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & x[54];
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & x[27];
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & ~x[17];
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & x[52];
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & ~x[14];
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & ~x[32];
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & x[54];
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & ~x[15];
			partial_clause[9][100] 	= partial_clause_prev[9][100] & ~x[51] & ~x[53];
			partial_clause[9][101] 	= partial_clause_prev[9][101] & 1'b1;
			partial_clause[9][102] 	= partial_clause_prev[9][102] & 1'b1;
			partial_clause[9][103] 	= partial_clause_prev[9][103] & 1'b1;
			partial_clause[9][104] 	= partial_clause_prev[9][104] & 1'b1;
			partial_clause[9][105] 	= partial_clause_prev[9][105] & 1'b1;
			partial_clause[9][106] 	= partial_clause_prev[9][106] & 1'b1;
			partial_clause[9][107] 	= partial_clause_prev[9][107] & 1'b1;
			partial_clause[9][108] 	= partial_clause_prev[9][108] & 1'b1;
			partial_clause[9][109] 	= partial_clause_prev[9][109] & 1'b1;
			partial_clause[9][110] 	= partial_clause_prev[9][110] & 1'b1;
			partial_clause[9][111] 	= partial_clause_prev[9][111] & 1'b1;
			partial_clause[9][112] 	= partial_clause_prev[9][112] & 1'b1;
			partial_clause[9][113] 	= partial_clause_prev[9][113] & 1'b1;
			partial_clause[9][114] 	= partial_clause_prev[9][114] & 1'b1;
			partial_clause[9][115] 	= partial_clause_prev[9][115] & 1'b1;
			partial_clause[9][116] 	= partial_clause_prev[9][116] & ~x[24];
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & 1'b1;
			partial_clause[9][119] 	= partial_clause_prev[9][119] & 1'b1;
			partial_clause[9][120] 	= partial_clause_prev[9][120] & 1'b1;
			partial_clause[9][121] 	= partial_clause_prev[9][121] & 1'b1;
			partial_clause[9][122] 	= partial_clause_prev[9][122] & 1'b1;
			partial_clause[9][123] 	= partial_clause_prev[9][123] & 1'b1;
			partial_clause[9][124] 	= partial_clause_prev[9][124] & ~x[39] & ~x[40];
			partial_clause[9][125] 	= partial_clause_prev[9][125] & 1'b1;
			partial_clause[9][126] 	= partial_clause_prev[9][126] & 1'b1;
			partial_clause[9][127] 	= partial_clause_prev[9][127] & 1'b1;
			partial_clause[9][128] 	= partial_clause_prev[9][128] & 1'b1;
			partial_clause[9][129] 	= partial_clause_prev[9][129] & 1'b1;
			partial_clause[9][130] 	= partial_clause_prev[9][130] & 1'b1;
			partial_clause[9][131] 	= partial_clause_prev[9][131] & 1'b1;
			partial_clause[9][132] 	= partial_clause_prev[9][132] & 1'b1;
			partial_clause[9][133] 	= partial_clause_prev[9][133] & 1'b1;
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & 1'b1;
			partial_clause[9][138] 	= partial_clause_prev[9][138] & 1'b1;
			partial_clause[9][139] 	= partial_clause_prev[9][139] & 1'b1;
			partial_clause[9][140] 	= partial_clause_prev[9][140] & 1'b1;
			partial_clause[9][141] 	= partial_clause_prev[9][141] & 1'b1;
			partial_clause[9][142] 	= partial_clause_prev[9][142] & 1'b1;
			partial_clause[9][143] 	= partial_clause_prev[9][143] & 1'b1;
			partial_clause[9][144] 	= partial_clause_prev[9][144] & 1'b1;
			partial_clause[9][145] 	= partial_clause_prev[9][145] & 1'b1;
			partial_clause[9][146] 	= partial_clause_prev[9][146] & 1'b1;
			partial_clause[9][147] 	= partial_clause_prev[9][147] & 1'b1;
			partial_clause[9][148] 	= partial_clause_prev[9][148] & 1'b1;
			partial_clause[9][149] 	= partial_clause_prev[9][149] & 1'b1;
			partial_clause[9][150] 	= partial_clause_prev[9][150] & 1'b1;
			partial_clause[9][151] 	= partial_clause_prev[9][151] & 1'b1;
			partial_clause[9][152] 	= partial_clause_prev[9][152] & 1'b1;
			partial_clause[9][153] 	= partial_clause_prev[9][153] & 1'b1;
			partial_clause[9][154] 	= partial_clause_prev[9][154] & 1'b1;
			partial_clause[9][155] 	= partial_clause_prev[9][155] & 1'b1;
			partial_clause[9][156] 	= partial_clause_prev[9][156] & 1'b1;
			partial_clause[9][157] 	= partial_clause_prev[9][157] & 1'b1;
			partial_clause[9][158] 	= partial_clause_prev[9][158] & 1'b1;
			partial_clause[9][159] 	= partial_clause_prev[9][159] & 1'b1;
			partial_clause[9][160] 	= partial_clause_prev[9][160] & 1'b1;
			partial_clause[9][161] 	= partial_clause_prev[9][161] & 1'b1;
			partial_clause[9][162] 	= partial_clause_prev[9][162] & 1'b1;
			partial_clause[9][163] 	= partial_clause_prev[9][163] & 1'b1;
			partial_clause[9][164] 	= partial_clause_prev[9][164] & 1'b1;
			partial_clause[9][165] 	= partial_clause_prev[9][165] & 1'b1;
			partial_clause[9][166] 	= partial_clause_prev[9][166] & 1'b1;
			partial_clause[9][167] 	= partial_clause_prev[9][167] & 1'b1;
			partial_clause[9][168] 	= partial_clause_prev[9][168] & ~x[39] & ~x[42];
			partial_clause[9][169] 	= partial_clause_prev[9][169] & 1'b1;
			partial_clause[9][170] 	= partial_clause_prev[9][170] & 1'b1;
			partial_clause[9][171] 	= partial_clause_prev[9][171] & 1'b1;
			partial_clause[9][172] 	= partial_clause_prev[9][172] & 1'b1;
			partial_clause[9][173] 	= partial_clause_prev[9][173] & 1'b1;
			partial_clause[9][174] 	= partial_clause_prev[9][174] & 1'b1;
			partial_clause[9][175] 	= partial_clause_prev[9][175] & 1'b1;
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & 1'b1;
			partial_clause[9][178] 	= partial_clause_prev[9][178] & 1'b1;
			partial_clause[9][179] 	= partial_clause_prev[9][179] & 1'b1;
			partial_clause[9][180] 	= partial_clause_prev[9][180] & 1'b1;
			partial_clause[9][181] 	= partial_clause_prev[9][181] & 1'b1;
			partial_clause[9][182] 	= partial_clause_prev[9][182] & 1'b1;
			partial_clause[9][183] 	= partial_clause_prev[9][183] & 1'b1;
			partial_clause[9][184] 	= partial_clause_prev[9][184] & 1'b1;
			partial_clause[9][185] 	= partial_clause_prev[9][185] & 1'b1;
			partial_clause[9][186] 	= partial_clause_prev[9][186] & 1'b1;
			partial_clause[9][187] 	= partial_clause_prev[9][187] & 1'b1;
			partial_clause[9][188] 	= partial_clause_prev[9][188] & 1'b1;
			partial_clause[9][189] 	= partial_clause_prev[9][189] & 1'b1;
			partial_clause[9][190] 	= partial_clause_prev[9][190] & 1'b1;
			partial_clause[9][191] 	= partial_clause_prev[9][191] & 1'b1;
			partial_clause[9][192] 	= partial_clause_prev[9][192] & 1'b1;
			partial_clause[9][193] 	= partial_clause_prev[9][193] & 1'b1;
			partial_clause[9][194] 	= partial_clause_prev[9][194] & 1'b1;
			partial_clause[9][195] 	= partial_clause_prev[9][195] & 1'b1;
			partial_clause[9][196] 	= partial_clause_prev[9][196] & ~x[53];
			partial_clause[9][197] 	= partial_clause_prev[9][197] & 1'b1;
			partial_clause[9][198] 	= partial_clause_prev[9][198] & 1'b1;
			partial_clause[9][199] 	= partial_clause_prev[9][199] & 1'b1;
		end
	end
endmodule


module HCB_11 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & ~x[8];
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & ~x[8];
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & x[60];
			partial_clause[0][20] 	= partial_clause_prev[0][20] & x[3];
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & ~x[8];
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & x[62];
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & ~x[12];
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & ~x[13];
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & ~x[6];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & x[43];
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			partial_clause[0][100] 	= partial_clause_prev[0][100] & 1'b1;
			partial_clause[0][101] 	= partial_clause_prev[0][101] & 1'b1;
			partial_clause[0][102] 	= partial_clause_prev[0][102] & 1'b1;
			partial_clause[0][103] 	= partial_clause_prev[0][103] & x[10];
			partial_clause[0][104] 	= partial_clause_prev[0][104] & 1'b1;
			partial_clause[0][105] 	= partial_clause_prev[0][105] & 1'b1;
			partial_clause[0][106] 	= partial_clause_prev[0][106] & 1'b1;
			partial_clause[0][107] 	= partial_clause_prev[0][107] & 1'b1;
			partial_clause[0][108] 	= partial_clause_prev[0][108] & 1'b1;
			partial_clause[0][109] 	= partial_clause_prev[0][109] & 1'b1;
			partial_clause[0][110] 	= partial_clause_prev[0][110] & ~x[22];
			partial_clause[0][111] 	= partial_clause_prev[0][111] & 1'b1;
			partial_clause[0][112] 	= partial_clause_prev[0][112] & 1'b1;
			partial_clause[0][113] 	= partial_clause_prev[0][113] & 1'b1;
			partial_clause[0][114] 	= partial_clause_prev[0][114] & 1'b1;
			partial_clause[0][115] 	= partial_clause_prev[0][115] & x[6];
			partial_clause[0][116] 	= partial_clause_prev[0][116] & 1'b1;
			partial_clause[0][117] 	= partial_clause_prev[0][117] & 1'b1;
			partial_clause[0][118] 	= partial_clause_prev[0][118] & 1'b1;
			partial_clause[0][119] 	= partial_clause_prev[0][119] & 1'b1;
			partial_clause[0][120] 	= partial_clause_prev[0][120] & 1'b1;
			partial_clause[0][121] 	= partial_clause_prev[0][121] & 1'b1;
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & 1'b1;
			partial_clause[0][124] 	= partial_clause_prev[0][124] & 1'b1;
			partial_clause[0][125] 	= partial_clause_prev[0][125] & 1'b1;
			partial_clause[0][126] 	= partial_clause_prev[0][126] & 1'b1;
			partial_clause[0][127] 	= partial_clause_prev[0][127] & 1'b1;
			partial_clause[0][128] 	= partial_clause_prev[0][128] & 1'b1;
			partial_clause[0][129] 	= partial_clause_prev[0][129] & 1'b1;
			partial_clause[0][130] 	= partial_clause_prev[0][130] & 1'b1;
			partial_clause[0][131] 	= partial_clause_prev[0][131] & 1'b1;
			partial_clause[0][132] 	= partial_clause_prev[0][132] & 1'b1;
			partial_clause[0][133] 	= partial_clause_prev[0][133] & x[11];
			partial_clause[0][134] 	= partial_clause_prev[0][134] & 1'b1;
			partial_clause[0][135] 	= partial_clause_prev[0][135] & 1'b1;
			partial_clause[0][136] 	= partial_clause_prev[0][136] & 1'b1;
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & 1'b1;
			partial_clause[0][139] 	= partial_clause_prev[0][139] & 1'b1;
			partial_clause[0][140] 	= partial_clause_prev[0][140] & 1'b1;
			partial_clause[0][141] 	= partial_clause_prev[0][141] & 1'b1;
			partial_clause[0][142] 	= partial_clause_prev[0][142] & 1'b1;
			partial_clause[0][143] 	= partial_clause_prev[0][143] & 1'b1;
			partial_clause[0][144] 	= partial_clause_prev[0][144] & 1'b1;
			partial_clause[0][145] 	= partial_clause_prev[0][145] & 1'b1;
			partial_clause[0][146] 	= partial_clause_prev[0][146] & 1'b1;
			partial_clause[0][147] 	= partial_clause_prev[0][147] & 1'b1;
			partial_clause[0][148] 	= partial_clause_prev[0][148] & 1'b1;
			partial_clause[0][149] 	= partial_clause_prev[0][149] & 1'b1;
			partial_clause[0][150] 	= partial_clause_prev[0][150] & 1'b1;
			partial_clause[0][151] 	= partial_clause_prev[0][151] & 1'b1;
			partial_clause[0][152] 	= partial_clause_prev[0][152] & 1'b1;
			partial_clause[0][153] 	= partial_clause_prev[0][153] & 1'b1;
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & 1'b1;
			partial_clause[0][156] 	= partial_clause_prev[0][156] & 1'b1;
			partial_clause[0][157] 	= partial_clause_prev[0][157] & 1'b1;
			partial_clause[0][158] 	= partial_clause_prev[0][158] & 1'b1;
			partial_clause[0][159] 	= partial_clause_prev[0][159] & 1'b1;
			partial_clause[0][160] 	= partial_clause_prev[0][160] & 1'b1;
			partial_clause[0][161] 	= partial_clause_prev[0][161] & 1'b1;
			partial_clause[0][162] 	= partial_clause_prev[0][162] & 1'b1;
			partial_clause[0][163] 	= partial_clause_prev[0][163] & x[10];
			partial_clause[0][164] 	= partial_clause_prev[0][164] & 1'b1;
			partial_clause[0][165] 	= partial_clause_prev[0][165] & 1'b1;
			partial_clause[0][166] 	= partial_clause_prev[0][166] & 1'b1;
			partial_clause[0][167] 	= partial_clause_prev[0][167] & 1'b1;
			partial_clause[0][168] 	= partial_clause_prev[0][168] & 1'b1;
			partial_clause[0][169] 	= partial_clause_prev[0][169] & 1'b1;
			partial_clause[0][170] 	= partial_clause_prev[0][170] & 1'b1;
			partial_clause[0][171] 	= partial_clause_prev[0][171] & 1'b1;
			partial_clause[0][172] 	= partial_clause_prev[0][172] & 1'b1;
			partial_clause[0][173] 	= partial_clause_prev[0][173] & 1'b1;
			partial_clause[0][174] 	= partial_clause_prev[0][174] & 1'b1;
			partial_clause[0][175] 	= partial_clause_prev[0][175] & x[7];
			partial_clause[0][176] 	= partial_clause_prev[0][176] & x[13];
			partial_clause[0][177] 	= partial_clause_prev[0][177] & 1'b1;
			partial_clause[0][178] 	= partial_clause_prev[0][178] & 1'b1;
			partial_clause[0][179] 	= partial_clause_prev[0][179] & 1'b1;
			partial_clause[0][180] 	= partial_clause_prev[0][180] & 1'b1;
			partial_clause[0][181] 	= partial_clause_prev[0][181] & x[8];
			partial_clause[0][182] 	= partial_clause_prev[0][182] & 1'b1;
			partial_clause[0][183] 	= partial_clause_prev[0][183] & 1'b1;
			partial_clause[0][184] 	= partial_clause_prev[0][184] & 1'b1;
			partial_clause[0][185] 	= partial_clause_prev[0][185] & 1'b1;
			partial_clause[0][186] 	= partial_clause_prev[0][186] & 1'b1;
			partial_clause[0][187] 	= partial_clause_prev[0][187] & 1'b1;
			partial_clause[0][188] 	= partial_clause_prev[0][188] & 1'b1;
			partial_clause[0][189] 	= partial_clause_prev[0][189] & 1'b1;
			partial_clause[0][190] 	= partial_clause_prev[0][190] & x[7];
			partial_clause[0][191] 	= partial_clause_prev[0][191] & 1'b1;
			partial_clause[0][192] 	= partial_clause_prev[0][192] & 1'b1;
			partial_clause[0][193] 	= partial_clause_prev[0][193] & 1'b1;
			partial_clause[0][194] 	= partial_clause_prev[0][194] & 1'b1;
			partial_clause[0][195] 	= partial_clause_prev[0][195] & 1'b1;
			partial_clause[0][196] 	= partial_clause_prev[0][196] & 1'b1;
			partial_clause[0][197] 	= partial_clause_prev[0][197] & 1'b1;
			partial_clause[0][198] 	= partial_clause_prev[0][198] & 1'b1;
			partial_clause[0][199] 	= partial_clause_prev[0][199] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & x[50];
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & x[24];
			partial_clause[1][12] 	= partial_clause_prev[1][12] & x[52];
			partial_clause[1][13] 	= partial_clause_prev[1][13] & x[17];
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & x[60];
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & x[1];
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & 1'b1;
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & x[19];
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & 1'b1;
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & x[48];
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & ~x[10];
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & x[28];
			partial_clause[1][92] 	= partial_clause_prev[1][92] & x[57];
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			partial_clause[1][100] 	= partial_clause_prev[1][100] & 1'b1;
			partial_clause[1][101] 	= partial_clause_prev[1][101] & 1'b1;
			partial_clause[1][102] 	= partial_clause_prev[1][102] & 1'b1;
			partial_clause[1][103] 	= partial_clause_prev[1][103] & 1'b1;
			partial_clause[1][104] 	= partial_clause_prev[1][104] & 1'b1;
			partial_clause[1][105] 	= partial_clause_prev[1][105] & 1'b1;
			partial_clause[1][106] 	= partial_clause_prev[1][106] & 1'b1;
			partial_clause[1][107] 	= partial_clause_prev[1][107] & 1'b1;
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & 1'b1;
			partial_clause[1][110] 	= partial_clause_prev[1][110] & 1'b1;
			partial_clause[1][111] 	= partial_clause_prev[1][111] & 1'b1;
			partial_clause[1][112] 	= partial_clause_prev[1][112] & 1'b1;
			partial_clause[1][113] 	= partial_clause_prev[1][113] & 1'b1;
			partial_clause[1][114] 	= partial_clause_prev[1][114] & 1'b1;
			partial_clause[1][115] 	= partial_clause_prev[1][115] & 1'b1;
			partial_clause[1][116] 	= partial_clause_prev[1][116] & 1'b1;
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & 1'b1;
			partial_clause[1][119] 	= partial_clause_prev[1][119] & 1'b1;
			partial_clause[1][120] 	= partial_clause_prev[1][120] & 1'b1;
			partial_clause[1][121] 	= partial_clause_prev[1][121] & 1'b1;
			partial_clause[1][122] 	= partial_clause_prev[1][122] & 1'b1;
			partial_clause[1][123] 	= partial_clause_prev[1][123] & 1'b1;
			partial_clause[1][124] 	= partial_clause_prev[1][124] & 1'b1;
			partial_clause[1][125] 	= partial_clause_prev[1][125] & 1'b1;
			partial_clause[1][126] 	= partial_clause_prev[1][126] & 1'b1;
			partial_clause[1][127] 	= partial_clause_prev[1][127] & 1'b1;
			partial_clause[1][128] 	= partial_clause_prev[1][128] & 1'b1;
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & 1'b1;
			partial_clause[1][131] 	= partial_clause_prev[1][131] & 1'b1;
			partial_clause[1][132] 	= partial_clause_prev[1][132] & 1'b1;
			partial_clause[1][133] 	= partial_clause_prev[1][133] & 1'b1;
			partial_clause[1][134] 	= partial_clause_prev[1][134] & 1'b1;
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & 1'b1;
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & 1'b1;
			partial_clause[1][139] 	= partial_clause_prev[1][139] & 1'b1;
			partial_clause[1][140] 	= partial_clause_prev[1][140] & x[6];
			partial_clause[1][141] 	= partial_clause_prev[1][141] & 1'b1;
			partial_clause[1][142] 	= partial_clause_prev[1][142] & 1'b1;
			partial_clause[1][143] 	= partial_clause_prev[1][143] & 1'b1;
			partial_clause[1][144] 	= partial_clause_prev[1][144] & 1'b1;
			partial_clause[1][145] 	= partial_clause_prev[1][145] & 1'b1;
			partial_clause[1][146] 	= partial_clause_prev[1][146] & 1'b1;
			partial_clause[1][147] 	= partial_clause_prev[1][147] & 1'b1;
			partial_clause[1][148] 	= partial_clause_prev[1][148] & 1'b1;
			partial_clause[1][149] 	= partial_clause_prev[1][149] & 1'b1;
			partial_clause[1][150] 	= partial_clause_prev[1][150] & ~x[1];
			partial_clause[1][151] 	= partial_clause_prev[1][151] & 1'b1;
			partial_clause[1][152] 	= partial_clause_prev[1][152] & 1'b1;
			partial_clause[1][153] 	= partial_clause_prev[1][153] & 1'b1;
			partial_clause[1][154] 	= partial_clause_prev[1][154] & 1'b1;
			partial_clause[1][155] 	= partial_clause_prev[1][155] & 1'b1;
			partial_clause[1][156] 	= partial_clause_prev[1][156] & 1'b1;
			partial_clause[1][157] 	= partial_clause_prev[1][157] & 1'b1;
			partial_clause[1][158] 	= partial_clause_prev[1][158] & 1'b1;
			partial_clause[1][159] 	= partial_clause_prev[1][159] & 1'b1;
			partial_clause[1][160] 	= partial_clause_prev[1][160] & 1'b1;
			partial_clause[1][161] 	= partial_clause_prev[1][161] & 1'b1;
			partial_clause[1][162] 	= partial_clause_prev[1][162] & 1'b1;
			partial_clause[1][163] 	= partial_clause_prev[1][163] & 1'b1;
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & 1'b1;
			partial_clause[1][166] 	= partial_clause_prev[1][166] & x[6];
			partial_clause[1][167] 	= partial_clause_prev[1][167] & 1'b1;
			partial_clause[1][168] 	= partial_clause_prev[1][168] & 1'b1;
			partial_clause[1][169] 	= partial_clause_prev[1][169] & 1'b1;
			partial_clause[1][170] 	= partial_clause_prev[1][170] & 1'b1;
			partial_clause[1][171] 	= partial_clause_prev[1][171] & 1'b1;
			partial_clause[1][172] 	= partial_clause_prev[1][172] & 1'b1;
			partial_clause[1][173] 	= partial_clause_prev[1][173] & 1'b1;
			partial_clause[1][174] 	= partial_clause_prev[1][174] & 1'b1;
			partial_clause[1][175] 	= partial_clause_prev[1][175] & 1'b1;
			partial_clause[1][176] 	= partial_clause_prev[1][176] & 1'b1;
			partial_clause[1][177] 	= partial_clause_prev[1][177] & 1'b1;
			partial_clause[1][178] 	= partial_clause_prev[1][178] & 1'b1;
			partial_clause[1][179] 	= partial_clause_prev[1][179] & 1'b1;
			partial_clause[1][180] 	= partial_clause_prev[1][180] & 1'b1;
			partial_clause[1][181] 	= partial_clause_prev[1][181] & 1'b1;
			partial_clause[1][182] 	= partial_clause_prev[1][182] & 1'b1;
			partial_clause[1][183] 	= partial_clause_prev[1][183] & 1'b1;
			partial_clause[1][184] 	= partial_clause_prev[1][184] & 1'b1;
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & 1'b1;
			partial_clause[1][187] 	= partial_clause_prev[1][187] & 1'b1;
			partial_clause[1][188] 	= partial_clause_prev[1][188] & 1'b1;
			partial_clause[1][189] 	= partial_clause_prev[1][189] & 1'b1;
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & 1'b1;
			partial_clause[1][192] 	= partial_clause_prev[1][192] & 1'b1;
			partial_clause[1][193] 	= partial_clause_prev[1][193] & 1'b1;
			partial_clause[1][194] 	= partial_clause_prev[1][194] & 1'b1;
			partial_clause[1][195] 	= partial_clause_prev[1][195] & 1'b1;
			partial_clause[1][196] 	= partial_clause_prev[1][196] & 1'b1;
			partial_clause[1][197] 	= partial_clause_prev[1][197] & 1'b1;
			partial_clause[1][198] 	= partial_clause_prev[1][198] & 1'b1;
			partial_clause[1][199] 	= partial_clause_prev[1][199] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & ~x[4];
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & ~x[6];
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & 1'b1;
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & ~x[3];
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			partial_clause[2][100] 	= partial_clause_prev[2][100] & 1'b1;
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & 1'b1;
			partial_clause[2][103] 	= partial_clause_prev[2][103] & 1'b1;
			partial_clause[2][104] 	= partial_clause_prev[2][104] & 1'b1;
			partial_clause[2][105] 	= partial_clause_prev[2][105] & 1'b1;
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & 1'b1;
			partial_clause[2][108] 	= partial_clause_prev[2][108] & 1'b1;
			partial_clause[2][109] 	= partial_clause_prev[2][109] & x[8];
			partial_clause[2][110] 	= partial_clause_prev[2][110] & 1'b1;
			partial_clause[2][111] 	= partial_clause_prev[2][111] & 1'b1;
			partial_clause[2][112] 	= partial_clause_prev[2][112] & 1'b1;
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & 1'b1;
			partial_clause[2][115] 	= partial_clause_prev[2][115] & 1'b1;
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & 1'b1;
			partial_clause[2][118] 	= partial_clause_prev[2][118] & 1'b1;
			partial_clause[2][119] 	= partial_clause_prev[2][119] & 1'b1;
			partial_clause[2][120] 	= partial_clause_prev[2][120] & 1'b1;
			partial_clause[2][121] 	= partial_clause_prev[2][121] & 1'b1;
			partial_clause[2][122] 	= partial_clause_prev[2][122] & 1'b1;
			partial_clause[2][123] 	= partial_clause_prev[2][123] & 1'b1;
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & 1'b1;
			partial_clause[2][126] 	= partial_clause_prev[2][126] & 1'b1;
			partial_clause[2][127] 	= partial_clause_prev[2][127] & 1'b1;
			partial_clause[2][128] 	= partial_clause_prev[2][128] & 1'b1;
			partial_clause[2][129] 	= partial_clause_prev[2][129] & x[10];
			partial_clause[2][130] 	= partial_clause_prev[2][130] & x[6];
			partial_clause[2][131] 	= partial_clause_prev[2][131] & 1'b1;
			partial_clause[2][132] 	= partial_clause_prev[2][132] & 1'b1;
			partial_clause[2][133] 	= partial_clause_prev[2][133] & x[5];
			partial_clause[2][134] 	= partial_clause_prev[2][134] & x[8];
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & 1'b1;
			partial_clause[2][137] 	= partial_clause_prev[2][137] & 1'b1;
			partial_clause[2][138] 	= partial_clause_prev[2][138] & 1'b1;
			partial_clause[2][139] 	= partial_clause_prev[2][139] & 1'b1;
			partial_clause[2][140] 	= partial_clause_prev[2][140] & 1'b1;
			partial_clause[2][141] 	= partial_clause_prev[2][141] & 1'b1;
			partial_clause[2][142] 	= partial_clause_prev[2][142] & 1'b1;
			partial_clause[2][143] 	= partial_clause_prev[2][143] & 1'b1;
			partial_clause[2][144] 	= partial_clause_prev[2][144] & 1'b1;
			partial_clause[2][145] 	= partial_clause_prev[2][145] & 1'b1;
			partial_clause[2][146] 	= partial_clause_prev[2][146] & 1'b1;
			partial_clause[2][147] 	= partial_clause_prev[2][147] & x[7];
			partial_clause[2][148] 	= partial_clause_prev[2][148] & 1'b1;
			partial_clause[2][149] 	= partial_clause_prev[2][149] & 1'b1;
			partial_clause[2][150] 	= partial_clause_prev[2][150] & 1'b1;
			partial_clause[2][151] 	= partial_clause_prev[2][151] & 1'b1;
			partial_clause[2][152] 	= partial_clause_prev[2][152] & 1'b1;
			partial_clause[2][153] 	= partial_clause_prev[2][153] & 1'b1;
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & 1'b1;
			partial_clause[2][156] 	= partial_clause_prev[2][156] & 1'b1;
			partial_clause[2][157] 	= partial_clause_prev[2][157] & 1'b1;
			partial_clause[2][158] 	= partial_clause_prev[2][158] & 1'b1;
			partial_clause[2][159] 	= partial_clause_prev[2][159] & 1'b1;
			partial_clause[2][160] 	= partial_clause_prev[2][160] & 1'b1;
			partial_clause[2][161] 	= partial_clause_prev[2][161] & 1'b1;
			partial_clause[2][162] 	= partial_clause_prev[2][162] & 1'b1;
			partial_clause[2][163] 	= partial_clause_prev[2][163] & 1'b1;
			partial_clause[2][164] 	= partial_clause_prev[2][164] & 1'b1;
			partial_clause[2][165] 	= partial_clause_prev[2][165] & 1'b1;
			partial_clause[2][166] 	= partial_clause_prev[2][166] & 1'b1;
			partial_clause[2][167] 	= partial_clause_prev[2][167] & 1'b1;
			partial_clause[2][168] 	= partial_clause_prev[2][168] & 1'b1;
			partial_clause[2][169] 	= partial_clause_prev[2][169] & 1'b1;
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & 1'b1;
			partial_clause[2][173] 	= partial_clause_prev[2][173] & 1'b1;
			partial_clause[2][174] 	= partial_clause_prev[2][174] & 1'b1;
			partial_clause[2][175] 	= partial_clause_prev[2][175] & 1'b1;
			partial_clause[2][176] 	= partial_clause_prev[2][176] & 1'b1;
			partial_clause[2][177] 	= partial_clause_prev[2][177] & 1'b1;
			partial_clause[2][178] 	= partial_clause_prev[2][178] & 1'b1;
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & x[4];
			partial_clause[2][181] 	= partial_clause_prev[2][181] & 1'b1;
			partial_clause[2][182] 	= partial_clause_prev[2][182] & 1'b1;
			partial_clause[2][183] 	= partial_clause_prev[2][183] & 1'b1;
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & x[4];
			partial_clause[2][186] 	= partial_clause_prev[2][186] & 1'b1;
			partial_clause[2][187] 	= partial_clause_prev[2][187] & 1'b1;
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & 1'b1;
			partial_clause[2][190] 	= partial_clause_prev[2][190] & 1'b1;
			partial_clause[2][191] 	= partial_clause_prev[2][191] & x[5];
			partial_clause[2][192] 	= partial_clause_prev[2][192] & 1'b1;
			partial_clause[2][193] 	= partial_clause_prev[2][193] & 1'b1;
			partial_clause[2][194] 	= partial_clause_prev[2][194] & 1'b1;
			partial_clause[2][195] 	= partial_clause_prev[2][195] & 1'b1;
			partial_clause[2][196] 	= partial_clause_prev[2][196] & 1'b1;
			partial_clause[2][197] 	= partial_clause_prev[2][197] & x[2];
			partial_clause[2][198] 	= partial_clause_prev[2][198] & 1'b1;
			partial_clause[2][199] 	= partial_clause_prev[2][199] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & x[1];
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & x[3];
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & x[6];
			partial_clause[3][21] 	= partial_clause_prev[3][21] & ~x[38];
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & x[0];
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[13];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & x[5];
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			partial_clause[3][100] 	= partial_clause_prev[3][100] & 1'b1;
			partial_clause[3][101] 	= partial_clause_prev[3][101] & 1'b1;
			partial_clause[3][102] 	= partial_clause_prev[3][102] & 1'b1;
			partial_clause[3][103] 	= partial_clause_prev[3][103] & 1'b1;
			partial_clause[3][104] 	= partial_clause_prev[3][104] & 1'b1;
			partial_clause[3][105] 	= partial_clause_prev[3][105] & 1'b1;
			partial_clause[3][106] 	= partial_clause_prev[3][106] & ~x[12];
			partial_clause[3][107] 	= partial_clause_prev[3][107] & 1'b1;
			partial_clause[3][108] 	= partial_clause_prev[3][108] & 1'b1;
			partial_clause[3][109] 	= partial_clause_prev[3][109] & 1'b1;
			partial_clause[3][110] 	= partial_clause_prev[3][110] & 1'b1;
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & 1'b1;
			partial_clause[3][113] 	= partial_clause_prev[3][113] & 1'b1;
			partial_clause[3][114] 	= partial_clause_prev[3][114] & 1'b1;
			partial_clause[3][115] 	= partial_clause_prev[3][115] & 1'b1;
			partial_clause[3][116] 	= partial_clause_prev[3][116] & 1'b1;
			partial_clause[3][117] 	= partial_clause_prev[3][117] & 1'b1;
			partial_clause[3][118] 	= partial_clause_prev[3][118] & 1'b1;
			partial_clause[3][119] 	= partial_clause_prev[3][119] & 1'b1;
			partial_clause[3][120] 	= partial_clause_prev[3][120] & 1'b1;
			partial_clause[3][121] 	= partial_clause_prev[3][121] & 1'b1;
			partial_clause[3][122] 	= partial_clause_prev[3][122] & 1'b1;
			partial_clause[3][123] 	= partial_clause_prev[3][123] & 1'b1;
			partial_clause[3][124] 	= partial_clause_prev[3][124] & 1'b1;
			partial_clause[3][125] 	= partial_clause_prev[3][125] & 1'b1;
			partial_clause[3][126] 	= partial_clause_prev[3][126] & 1'b1;
			partial_clause[3][127] 	= partial_clause_prev[3][127] & 1'b1;
			partial_clause[3][128] 	= partial_clause_prev[3][128] & 1'b1;
			partial_clause[3][129] 	= partial_clause_prev[3][129] & x[46];
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & 1'b1;
			partial_clause[3][132] 	= partial_clause_prev[3][132] & 1'b1;
			partial_clause[3][133] 	= partial_clause_prev[3][133] & 1'b1;
			partial_clause[3][134] 	= partial_clause_prev[3][134] & 1'b1;
			partial_clause[3][135] 	= partial_clause_prev[3][135] & 1'b1;
			partial_clause[3][136] 	= partial_clause_prev[3][136] & 1'b1;
			partial_clause[3][137] 	= partial_clause_prev[3][137] & 1'b1;
			partial_clause[3][138] 	= partial_clause_prev[3][138] & 1'b1;
			partial_clause[3][139] 	= partial_clause_prev[3][139] & 1'b1;
			partial_clause[3][140] 	= partial_clause_prev[3][140] & 1'b1;
			partial_clause[3][141] 	= partial_clause_prev[3][141] & 1'b1;
			partial_clause[3][142] 	= partial_clause_prev[3][142] & 1'b1;
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & 1'b1;
			partial_clause[3][145] 	= partial_clause_prev[3][145] & 1'b1;
			partial_clause[3][146] 	= partial_clause_prev[3][146] & 1'b1;
			partial_clause[3][147] 	= partial_clause_prev[3][147] & 1'b1;
			partial_clause[3][148] 	= partial_clause_prev[3][148] & 1'b1;
			partial_clause[3][149] 	= partial_clause_prev[3][149] & 1'b1;
			partial_clause[3][150] 	= partial_clause_prev[3][150] & 1'b1;
			partial_clause[3][151] 	= partial_clause_prev[3][151] & ~x[8];
			partial_clause[3][152] 	= partial_clause_prev[3][152] & 1'b1;
			partial_clause[3][153] 	= partial_clause_prev[3][153] & x[39];
			partial_clause[3][154] 	= partial_clause_prev[3][154] & 1'b1;
			partial_clause[3][155] 	= partial_clause_prev[3][155] & 1'b1;
			partial_clause[3][156] 	= partial_clause_prev[3][156] & 1'b1;
			partial_clause[3][157] 	= partial_clause_prev[3][157] & 1'b1;
			partial_clause[3][158] 	= partial_clause_prev[3][158] & 1'b1;
			partial_clause[3][159] 	= partial_clause_prev[3][159] & 1'b1;
			partial_clause[3][160] 	= partial_clause_prev[3][160] & 1'b1;
			partial_clause[3][161] 	= partial_clause_prev[3][161] & x[14];
			partial_clause[3][162] 	= partial_clause_prev[3][162] & 1'b1;
			partial_clause[3][163] 	= partial_clause_prev[3][163] & 1'b1;
			partial_clause[3][164] 	= partial_clause_prev[3][164] & 1'b1;
			partial_clause[3][165] 	= partial_clause_prev[3][165] & 1'b1;
			partial_clause[3][166] 	= partial_clause_prev[3][166] & 1'b1;
			partial_clause[3][167] 	= partial_clause_prev[3][167] & 1'b1;
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & 1'b1;
			partial_clause[3][170] 	= partial_clause_prev[3][170] & 1'b1;
			partial_clause[3][171] 	= partial_clause_prev[3][171] & 1'b1;
			partial_clause[3][172] 	= partial_clause_prev[3][172] & 1'b1;
			partial_clause[3][173] 	= partial_clause_prev[3][173] & 1'b1;
			partial_clause[3][174] 	= partial_clause_prev[3][174] & 1'b1;
			partial_clause[3][175] 	= partial_clause_prev[3][175] & 1'b1;
			partial_clause[3][176] 	= partial_clause_prev[3][176] & 1'b1;
			partial_clause[3][177] 	= partial_clause_prev[3][177] & 1'b1;
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & 1'b1;
			partial_clause[3][180] 	= partial_clause_prev[3][180] & 1'b1;
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & 1'b1;
			partial_clause[3][183] 	= partial_clause_prev[3][183] & 1'b1;
			partial_clause[3][184] 	= partial_clause_prev[3][184] & 1'b1;
			partial_clause[3][185] 	= partial_clause_prev[3][185] & 1'b1;
			partial_clause[3][186] 	= partial_clause_prev[3][186] & 1'b1;
			partial_clause[3][187] 	= partial_clause_prev[3][187] & 1'b1;
			partial_clause[3][188] 	= partial_clause_prev[3][188] & 1'b1;
			partial_clause[3][189] 	= partial_clause_prev[3][189] & 1'b1;
			partial_clause[3][190] 	= partial_clause_prev[3][190] & 1'b1;
			partial_clause[3][191] 	= partial_clause_prev[3][191] & 1'b1;
			partial_clause[3][192] 	= partial_clause_prev[3][192] & 1'b1;
			partial_clause[3][193] 	= partial_clause_prev[3][193] & 1'b1;
			partial_clause[3][194] 	= partial_clause_prev[3][194] & 1'b1;
			partial_clause[3][195] 	= partial_clause_prev[3][195] & 1'b1;
			partial_clause[3][196] 	= partial_clause_prev[3][196] & x[20];
			partial_clause[3][197] 	= partial_clause_prev[3][197] & 1'b1;
			partial_clause[3][198] 	= partial_clause_prev[3][198] & 1'b1;
			partial_clause[3][199] 	= partial_clause_prev[3][199] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & ~x[7] & ~x[12];
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & ~x[10] & ~x[11];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & 1'b1;
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & x[23];
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & x[26];
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & 1'b1;
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & ~x[5];
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & ~x[10] & ~x[36];
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & x[22];
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & ~x[7] & ~x[8] & ~x[9];
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & ~x[38];
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & x[23];
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & ~x[6];
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			partial_clause[4][100] 	= partial_clause_prev[4][100] & 1'b1;
			partial_clause[4][101] 	= partial_clause_prev[4][101] & 1'b1;
			partial_clause[4][102] 	= partial_clause_prev[4][102] & 1'b1;
			partial_clause[4][103] 	= partial_clause_prev[4][103] & 1'b1;
			partial_clause[4][104] 	= partial_clause_prev[4][104] & 1'b1;
			partial_clause[4][105] 	= partial_clause_prev[4][105] & 1'b1;
			partial_clause[4][106] 	= partial_clause_prev[4][106] & 1'b1;
			partial_clause[4][107] 	= partial_clause_prev[4][107] & 1'b1;
			partial_clause[4][108] 	= partial_clause_prev[4][108] & 1'b1;
			partial_clause[4][109] 	= partial_clause_prev[4][109] & 1'b1;
			partial_clause[4][110] 	= partial_clause_prev[4][110] & 1'b1;
			partial_clause[4][111] 	= partial_clause_prev[4][111] & 1'b1;
			partial_clause[4][112] 	= partial_clause_prev[4][112] & 1'b1;
			partial_clause[4][113] 	= partial_clause_prev[4][113] & 1'b1;
			partial_clause[4][114] 	= partial_clause_prev[4][114] & 1'b1;
			partial_clause[4][115] 	= partial_clause_prev[4][115] & 1'b1;
			partial_clause[4][116] 	= partial_clause_prev[4][116] & 1'b1;
			partial_clause[4][117] 	= partial_clause_prev[4][117] & ~x[51];
			partial_clause[4][118] 	= partial_clause_prev[4][118] & 1'b1;
			partial_clause[4][119] 	= partial_clause_prev[4][119] & 1'b1;
			partial_clause[4][120] 	= partial_clause_prev[4][120] & 1'b1;
			partial_clause[4][121] 	= partial_clause_prev[4][121] & 1'b1;
			partial_clause[4][122] 	= partial_clause_prev[4][122] & 1'b1;
			partial_clause[4][123] 	= partial_clause_prev[4][123] & 1'b1;
			partial_clause[4][124] 	= partial_clause_prev[4][124] & x[38];
			partial_clause[4][125] 	= partial_clause_prev[4][125] & 1'b1;
			partial_clause[4][126] 	= partial_clause_prev[4][126] & x[13];
			partial_clause[4][127] 	= partial_clause_prev[4][127] & 1'b1;
			partial_clause[4][128] 	= partial_clause_prev[4][128] & 1'b1;
			partial_clause[4][129] 	= partial_clause_prev[4][129] & 1'b1;
			partial_clause[4][130] 	= partial_clause_prev[4][130] & 1'b1;
			partial_clause[4][131] 	= partial_clause_prev[4][131] & 1'b1;
			partial_clause[4][132] 	= partial_clause_prev[4][132] & 1'b1;
			partial_clause[4][133] 	= partial_clause_prev[4][133] & 1'b1;
			partial_clause[4][134] 	= partial_clause_prev[4][134] & x[35];
			partial_clause[4][135] 	= partial_clause_prev[4][135] & 1'b1;
			partial_clause[4][136] 	= partial_clause_prev[4][136] & 1'b1;
			partial_clause[4][137] 	= partial_clause_prev[4][137] & 1'b1;
			partial_clause[4][138] 	= partial_clause_prev[4][138] & 1'b1;
			partial_clause[4][139] 	= partial_clause_prev[4][139] & x[33];
			partial_clause[4][140] 	= partial_clause_prev[4][140] & 1'b1;
			partial_clause[4][141] 	= partial_clause_prev[4][141] & 1'b1;
			partial_clause[4][142] 	= partial_clause_prev[4][142] & 1'b1;
			partial_clause[4][143] 	= partial_clause_prev[4][143] & 1'b1;
			partial_clause[4][144] 	= partial_clause_prev[4][144] & 1'b1;
			partial_clause[4][145] 	= partial_clause_prev[4][145] & x[12];
			partial_clause[4][146] 	= partial_clause_prev[4][146] & 1'b1;
			partial_clause[4][147] 	= partial_clause_prev[4][147] & x[8];
			partial_clause[4][148] 	= partial_clause_prev[4][148] & 1'b1;
			partial_clause[4][149] 	= partial_clause_prev[4][149] & 1'b1;
			partial_clause[4][150] 	= partial_clause_prev[4][150] & 1'b1;
			partial_clause[4][151] 	= partial_clause_prev[4][151] & 1'b1;
			partial_clause[4][152] 	= partial_clause_prev[4][152] & 1'b1;
			partial_clause[4][153] 	= partial_clause_prev[4][153] & 1'b1;
			partial_clause[4][154] 	= partial_clause_prev[4][154] & 1'b1;
			partial_clause[4][155] 	= partial_clause_prev[4][155] & 1'b1;
			partial_clause[4][156] 	= partial_clause_prev[4][156] & 1'b1;
			partial_clause[4][157] 	= partial_clause_prev[4][157] & 1'b1;
			partial_clause[4][158] 	= partial_clause_prev[4][158] & 1'b1;
			partial_clause[4][159] 	= partial_clause_prev[4][159] & 1'b1;
			partial_clause[4][160] 	= partial_clause_prev[4][160] & 1'b1;
			partial_clause[4][161] 	= partial_clause_prev[4][161] & 1'b1;
			partial_clause[4][162] 	= partial_clause_prev[4][162] & 1'b1;
			partial_clause[4][163] 	= partial_clause_prev[4][163] & 1'b1;
			partial_clause[4][164] 	= partial_clause_prev[4][164] & 1'b1;
			partial_clause[4][165] 	= partial_clause_prev[4][165] & 1'b1;
			partial_clause[4][166] 	= partial_clause_prev[4][166] & 1'b1;
			partial_clause[4][167] 	= partial_clause_prev[4][167] & 1'b1;
			partial_clause[4][168] 	= partial_clause_prev[4][168] & x[12];
			partial_clause[4][169] 	= partial_clause_prev[4][169] & 1'b1;
			partial_clause[4][170] 	= partial_clause_prev[4][170] & 1'b1;
			partial_clause[4][171] 	= partial_clause_prev[4][171] & 1'b1;
			partial_clause[4][172] 	= partial_clause_prev[4][172] & 1'b1;
			partial_clause[4][173] 	= partial_clause_prev[4][173] & 1'b1;
			partial_clause[4][174] 	= partial_clause_prev[4][174] & 1'b1;
			partial_clause[4][175] 	= partial_clause_prev[4][175] & 1'b1;
			partial_clause[4][176] 	= partial_clause_prev[4][176] & x[8];
			partial_clause[4][177] 	= partial_clause_prev[4][177] & 1'b1;
			partial_clause[4][178] 	= partial_clause_prev[4][178] & 1'b1;
			partial_clause[4][179] 	= partial_clause_prev[4][179] & 1'b1;
			partial_clause[4][180] 	= partial_clause_prev[4][180] & 1'b1;
			partial_clause[4][181] 	= partial_clause_prev[4][181] & 1'b1;
			partial_clause[4][182] 	= partial_clause_prev[4][182] & 1'b1;
			partial_clause[4][183] 	= partial_clause_prev[4][183] & 1'b1;
			partial_clause[4][184] 	= partial_clause_prev[4][184] & 1'b1;
			partial_clause[4][185] 	= partial_clause_prev[4][185] & 1'b1;
			partial_clause[4][186] 	= partial_clause_prev[4][186] & 1'b1;
			partial_clause[4][187] 	= partial_clause_prev[4][187] & 1'b1;
			partial_clause[4][188] 	= partial_clause_prev[4][188] & 1'b1;
			partial_clause[4][189] 	= partial_clause_prev[4][189] & 1'b1;
			partial_clause[4][190] 	= partial_clause_prev[4][190] & 1'b1;
			partial_clause[4][191] 	= partial_clause_prev[4][191] & 1'b1;
			partial_clause[4][192] 	= partial_clause_prev[4][192] & 1'b1;
			partial_clause[4][193] 	= partial_clause_prev[4][193] & 1'b1;
			partial_clause[4][194] 	= partial_clause_prev[4][194] & 1'b1;
			partial_clause[4][195] 	= partial_clause_prev[4][195] & 1'b1;
			partial_clause[4][196] 	= partial_clause_prev[4][196] & 1'b1;
			partial_clause[4][197] 	= partial_clause_prev[4][197] & 1'b1;
			partial_clause[4][198] 	= partial_clause_prev[4][198] & 1'b1;
			partial_clause[4][199] 	= partial_clause_prev[4][199] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & ~x[47];
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & x[53];
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			partial_clause[5][100] 	= partial_clause_prev[5][100] & 1'b1;
			partial_clause[5][101] 	= partial_clause_prev[5][101] & x[34];
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & 1'b1;
			partial_clause[5][104] 	= partial_clause_prev[5][104] & 1'b1;
			partial_clause[5][105] 	= partial_clause_prev[5][105] & 1'b1;
			partial_clause[5][106] 	= partial_clause_prev[5][106] & 1'b1;
			partial_clause[5][107] 	= partial_clause_prev[5][107] & 1'b1;
			partial_clause[5][108] 	= partial_clause_prev[5][108] & 1'b1;
			partial_clause[5][109] 	= partial_clause_prev[5][109] & 1'b1;
			partial_clause[5][110] 	= partial_clause_prev[5][110] & 1'b1;
			partial_clause[5][111] 	= partial_clause_prev[5][111] & 1'b1;
			partial_clause[5][112] 	= partial_clause_prev[5][112] & 1'b1;
			partial_clause[5][113] 	= partial_clause_prev[5][113] & 1'b1;
			partial_clause[5][114] 	= partial_clause_prev[5][114] & 1'b1;
			partial_clause[5][115] 	= partial_clause_prev[5][115] & 1'b1;
			partial_clause[5][116] 	= partial_clause_prev[5][116] & x[39];
			partial_clause[5][117] 	= partial_clause_prev[5][117] & 1'b1;
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & 1'b1;
			partial_clause[5][120] 	= partial_clause_prev[5][120] & 1'b1;
			partial_clause[5][121] 	= partial_clause_prev[5][121] & 1'b1;
			partial_clause[5][122] 	= partial_clause_prev[5][122] & 1'b1;
			partial_clause[5][123] 	= partial_clause_prev[5][123] & 1'b1;
			partial_clause[5][124] 	= partial_clause_prev[5][124] & x[55];
			partial_clause[5][125] 	= partial_clause_prev[5][125] & 1'b1;
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & 1'b1;
			partial_clause[5][128] 	= partial_clause_prev[5][128] & 1'b1;
			partial_clause[5][129] 	= partial_clause_prev[5][129] & 1'b1;
			partial_clause[5][130] 	= partial_clause_prev[5][130] & 1'b1;
			partial_clause[5][131] 	= partial_clause_prev[5][131] & 1'b1;
			partial_clause[5][132] 	= partial_clause_prev[5][132] & 1'b1;
			partial_clause[5][133] 	= partial_clause_prev[5][133] & 1'b1;
			partial_clause[5][134] 	= partial_clause_prev[5][134] & 1'b1;
			partial_clause[5][135] 	= partial_clause_prev[5][135] & 1'b1;
			partial_clause[5][136] 	= partial_clause_prev[5][136] & 1'b1;
			partial_clause[5][137] 	= partial_clause_prev[5][137] & 1'b1;
			partial_clause[5][138] 	= partial_clause_prev[5][138] & 1'b1;
			partial_clause[5][139] 	= partial_clause_prev[5][139] & 1'b1;
			partial_clause[5][140] 	= partial_clause_prev[5][140] & 1'b1;
			partial_clause[5][141] 	= partial_clause_prev[5][141] & 1'b1;
			partial_clause[5][142] 	= partial_clause_prev[5][142] & 1'b1;
			partial_clause[5][143] 	= partial_clause_prev[5][143] & 1'b1;
			partial_clause[5][144] 	= partial_clause_prev[5][144] & 1'b1;
			partial_clause[5][145] 	= partial_clause_prev[5][145] & 1'b1;
			partial_clause[5][146] 	= partial_clause_prev[5][146] & 1'b1;
			partial_clause[5][147] 	= partial_clause_prev[5][147] & 1'b1;
			partial_clause[5][148] 	= partial_clause_prev[5][148] & 1'b1;
			partial_clause[5][149] 	= partial_clause_prev[5][149] & 1'b1;
			partial_clause[5][150] 	= partial_clause_prev[5][150] & 1'b1;
			partial_clause[5][151] 	= partial_clause_prev[5][151] & 1'b1;
			partial_clause[5][152] 	= partial_clause_prev[5][152] & 1'b1;
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & 1'b1;
			partial_clause[5][155] 	= partial_clause_prev[5][155] & 1'b1;
			partial_clause[5][156] 	= partial_clause_prev[5][156] & 1'b1;
			partial_clause[5][157] 	= partial_clause_prev[5][157] & 1'b1;
			partial_clause[5][158] 	= partial_clause_prev[5][158] & 1'b1;
			partial_clause[5][159] 	= partial_clause_prev[5][159] & 1'b1;
			partial_clause[5][160] 	= partial_clause_prev[5][160] & x[31];
			partial_clause[5][161] 	= partial_clause_prev[5][161] & 1'b1;
			partial_clause[5][162] 	= partial_clause_prev[5][162] & 1'b1;
			partial_clause[5][163] 	= partial_clause_prev[5][163] & 1'b1;
			partial_clause[5][164] 	= partial_clause_prev[5][164] & 1'b1;
			partial_clause[5][165] 	= partial_clause_prev[5][165] & 1'b1;
			partial_clause[5][166] 	= partial_clause_prev[5][166] & 1'b1;
			partial_clause[5][167] 	= partial_clause_prev[5][167] & 1'b1;
			partial_clause[5][168] 	= partial_clause_prev[5][168] & 1'b1;
			partial_clause[5][169] 	= partial_clause_prev[5][169] & 1'b1;
			partial_clause[5][170] 	= partial_clause_prev[5][170] & 1'b1;
			partial_clause[5][171] 	= partial_clause_prev[5][171] & 1'b1;
			partial_clause[5][172] 	= partial_clause_prev[5][172] & 1'b1;
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & 1'b1;
			partial_clause[5][175] 	= partial_clause_prev[5][175] & 1'b1;
			partial_clause[5][176] 	= partial_clause_prev[5][176] & 1'b1;
			partial_clause[5][177] 	= partial_clause_prev[5][177] & 1'b1;
			partial_clause[5][178] 	= partial_clause_prev[5][178] & 1'b1;
			partial_clause[5][179] 	= partial_clause_prev[5][179] & 1'b1;
			partial_clause[5][180] 	= partial_clause_prev[5][180] & 1'b1;
			partial_clause[5][181] 	= partial_clause_prev[5][181] & 1'b1;
			partial_clause[5][182] 	= partial_clause_prev[5][182] & 1'b1;
			partial_clause[5][183] 	= partial_clause_prev[5][183] & 1'b1;
			partial_clause[5][184] 	= partial_clause_prev[5][184] & 1'b1;
			partial_clause[5][185] 	= partial_clause_prev[5][185] & 1'b1;
			partial_clause[5][186] 	= partial_clause_prev[5][186] & 1'b1;
			partial_clause[5][187] 	= partial_clause_prev[5][187] & 1'b1;
			partial_clause[5][188] 	= partial_clause_prev[5][188] & 1'b1;
			partial_clause[5][189] 	= partial_clause_prev[5][189] & 1'b1;
			partial_clause[5][190] 	= partial_clause_prev[5][190] & 1'b1;
			partial_clause[5][191] 	= partial_clause_prev[5][191] & 1'b1;
			partial_clause[5][192] 	= partial_clause_prev[5][192] & 1'b1;
			partial_clause[5][193] 	= partial_clause_prev[5][193] & 1'b1;
			partial_clause[5][194] 	= partial_clause_prev[5][194] & 1'b1;
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & 1'b1;
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & 1'b1;
			partial_clause[5][199] 	= partial_clause_prev[5][199] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & x[3];
			partial_clause[6][16] 	= partial_clause_prev[6][16] & x[42];
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & ~x[44];
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & x[21];
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & x[21];
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			partial_clause[6][100] 	= partial_clause_prev[6][100] & 1'b1;
			partial_clause[6][101] 	= partial_clause_prev[6][101] & 1'b1;
			partial_clause[6][102] 	= partial_clause_prev[6][102] & 1'b1;
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & 1'b1;
			partial_clause[6][105] 	= partial_clause_prev[6][105] & 1'b1;
			partial_clause[6][106] 	= partial_clause_prev[6][106] & 1'b1;
			partial_clause[6][107] 	= partial_clause_prev[6][107] & 1'b1;
			partial_clause[6][108] 	= partial_clause_prev[6][108] & 1'b1;
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & 1'b1;
			partial_clause[6][111] 	= partial_clause_prev[6][111] & 1'b1;
			partial_clause[6][112] 	= partial_clause_prev[6][112] & 1'b1;
			partial_clause[6][113] 	= partial_clause_prev[6][113] & 1'b1;
			partial_clause[6][114] 	= partial_clause_prev[6][114] & 1'b1;
			partial_clause[6][115] 	= partial_clause_prev[6][115] & 1'b1;
			partial_clause[6][116] 	= partial_clause_prev[6][116] & 1'b1;
			partial_clause[6][117] 	= partial_clause_prev[6][117] & 1'b1;
			partial_clause[6][118] 	= partial_clause_prev[6][118] & 1'b1;
			partial_clause[6][119] 	= partial_clause_prev[6][119] & 1'b1;
			partial_clause[6][120] 	= partial_clause_prev[6][120] & 1'b1;
			partial_clause[6][121] 	= partial_clause_prev[6][121] & 1'b1;
			partial_clause[6][122] 	= partial_clause_prev[6][122] & 1'b1;
			partial_clause[6][123] 	= partial_clause_prev[6][123] & 1'b1;
			partial_clause[6][124] 	= partial_clause_prev[6][124] & 1'b1;
			partial_clause[6][125] 	= partial_clause_prev[6][125] & 1'b1;
			partial_clause[6][126] 	= partial_clause_prev[6][126] & 1'b1;
			partial_clause[6][127] 	= partial_clause_prev[6][127] & 1'b1;
			partial_clause[6][128] 	= partial_clause_prev[6][128] & 1'b1;
			partial_clause[6][129] 	= partial_clause_prev[6][129] & 1'b1;
			partial_clause[6][130] 	= partial_clause_prev[6][130] & 1'b1;
			partial_clause[6][131] 	= partial_clause_prev[6][131] & 1'b1;
			partial_clause[6][132] 	= partial_clause_prev[6][132] & 1'b1;
			partial_clause[6][133] 	= partial_clause_prev[6][133] & 1'b1;
			partial_clause[6][134] 	= partial_clause_prev[6][134] & 1'b1;
			partial_clause[6][135] 	= partial_clause_prev[6][135] & 1'b1;
			partial_clause[6][136] 	= partial_clause_prev[6][136] & ~x[48];
			partial_clause[6][137] 	= partial_clause_prev[6][137] & 1'b1;
			partial_clause[6][138] 	= partial_clause_prev[6][138] & 1'b1;
			partial_clause[6][139] 	= partial_clause_prev[6][139] & 1'b1;
			partial_clause[6][140] 	= partial_clause_prev[6][140] & 1'b1;
			partial_clause[6][141] 	= partial_clause_prev[6][141] & 1'b1;
			partial_clause[6][142] 	= partial_clause_prev[6][142] & 1'b1;
			partial_clause[6][143] 	= partial_clause_prev[6][143] & 1'b1;
			partial_clause[6][144] 	= partial_clause_prev[6][144] & 1'b1;
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & 1'b1;
			partial_clause[6][147] 	= partial_clause_prev[6][147] & 1'b1;
			partial_clause[6][148] 	= partial_clause_prev[6][148] & 1'b1;
			partial_clause[6][149] 	= partial_clause_prev[6][149] & 1'b1;
			partial_clause[6][150] 	= partial_clause_prev[6][150] & 1'b1;
			partial_clause[6][151] 	= partial_clause_prev[6][151] & 1'b1;
			partial_clause[6][152] 	= partial_clause_prev[6][152] & 1'b1;
			partial_clause[6][153] 	= partial_clause_prev[6][153] & ~x[29];
			partial_clause[6][154] 	= partial_clause_prev[6][154] & 1'b1;
			partial_clause[6][155] 	= partial_clause_prev[6][155] & 1'b1;
			partial_clause[6][156] 	= partial_clause_prev[6][156] & 1'b1;
			partial_clause[6][157] 	= partial_clause_prev[6][157] & 1'b1;
			partial_clause[6][158] 	= partial_clause_prev[6][158] & 1'b1;
			partial_clause[6][159] 	= partial_clause_prev[6][159] & 1'b1;
			partial_clause[6][160] 	= partial_clause_prev[6][160] & 1'b1;
			partial_clause[6][161] 	= partial_clause_prev[6][161] & 1'b1;
			partial_clause[6][162] 	= partial_clause_prev[6][162] & 1'b1;
			partial_clause[6][163] 	= partial_clause_prev[6][163] & 1'b1;
			partial_clause[6][164] 	= partial_clause_prev[6][164] & 1'b1;
			partial_clause[6][165] 	= partial_clause_prev[6][165] & 1'b1;
			partial_clause[6][166] 	= partial_clause_prev[6][166] & 1'b1;
			partial_clause[6][167] 	= partial_clause_prev[6][167] & 1'b1;
			partial_clause[6][168] 	= partial_clause_prev[6][168] & 1'b1;
			partial_clause[6][169] 	= partial_clause_prev[6][169] & 1'b1;
			partial_clause[6][170] 	= partial_clause_prev[6][170] & 1'b1;
			partial_clause[6][171] 	= partial_clause_prev[6][171] & 1'b1;
			partial_clause[6][172] 	= partial_clause_prev[6][172] & ~x[20];
			partial_clause[6][173] 	= partial_clause_prev[6][173] & 1'b1;
			partial_clause[6][174] 	= partial_clause_prev[6][174] & 1'b1;
			partial_clause[6][175] 	= partial_clause_prev[6][175] & 1'b1;
			partial_clause[6][176] 	= partial_clause_prev[6][176] & 1'b1;
			partial_clause[6][177] 	= partial_clause_prev[6][177] & 1'b1;
			partial_clause[6][178] 	= partial_clause_prev[6][178] & 1'b1;
			partial_clause[6][179] 	= partial_clause_prev[6][179] & 1'b1;
			partial_clause[6][180] 	= partial_clause_prev[6][180] & 1'b1;
			partial_clause[6][181] 	= partial_clause_prev[6][181] & 1'b1;
			partial_clause[6][182] 	= partial_clause_prev[6][182] & 1'b1;
			partial_clause[6][183] 	= partial_clause_prev[6][183] & 1'b1;
			partial_clause[6][184] 	= partial_clause_prev[6][184] & 1'b1;
			partial_clause[6][185] 	= partial_clause_prev[6][185] & 1'b1;
			partial_clause[6][186] 	= partial_clause_prev[6][186] & 1'b1;
			partial_clause[6][187] 	= partial_clause_prev[6][187] & 1'b1;
			partial_clause[6][188] 	= partial_clause_prev[6][188] & 1'b1;
			partial_clause[6][189] 	= partial_clause_prev[6][189] & 1'b1;
			partial_clause[6][190] 	= partial_clause_prev[6][190] & 1'b1;
			partial_clause[6][191] 	= partial_clause_prev[6][191] & 1'b1;
			partial_clause[6][192] 	= partial_clause_prev[6][192] & 1'b1;
			partial_clause[6][193] 	= partial_clause_prev[6][193] & 1'b1;
			partial_clause[6][194] 	= partial_clause_prev[6][194] & 1'b1;
			partial_clause[6][195] 	= partial_clause_prev[6][195] & 1'b1;
			partial_clause[6][196] 	= partial_clause_prev[6][196] & 1'b1;
			partial_clause[6][197] 	= partial_clause_prev[6][197] & 1'b1;
			partial_clause[6][198] 	= partial_clause_prev[6][198] & 1'b1;
			partial_clause[6][199] 	= partial_clause_prev[6][199] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & x[33];
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & x[8];
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & x[46];
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & x[59];
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & x[35];
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & x[13];
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & x[41];
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & x[10];
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & x[1];
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & x[33];
			partial_clause[7][61] 	= partial_clause_prev[7][61] & x[6];
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & x[11];
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & x[1];
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & x[37];
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & x[3];
			partial_clause[7][91] 	= partial_clause_prev[7][91] & x[26];
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & x[39];
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			partial_clause[7][100] 	= partial_clause_prev[7][100] & 1'b1;
			partial_clause[7][101] 	= partial_clause_prev[7][101] & 1'b1;
			partial_clause[7][102] 	= partial_clause_prev[7][102] & 1'b1;
			partial_clause[7][103] 	= partial_clause_prev[7][103] & 1'b1;
			partial_clause[7][104] 	= partial_clause_prev[7][104] & 1'b1;
			partial_clause[7][105] 	= partial_clause_prev[7][105] & 1'b1;
			partial_clause[7][106] 	= partial_clause_prev[7][106] & 1'b1;
			partial_clause[7][107] 	= partial_clause_prev[7][107] & 1'b1;
			partial_clause[7][108] 	= partial_clause_prev[7][108] & 1'b1;
			partial_clause[7][109] 	= partial_clause_prev[7][109] & 1'b1;
			partial_clause[7][110] 	= partial_clause_prev[7][110] & 1'b1;
			partial_clause[7][111] 	= partial_clause_prev[7][111] & 1'b1;
			partial_clause[7][112] 	= partial_clause_prev[7][112] & 1'b1;
			partial_clause[7][113] 	= partial_clause_prev[7][113] & 1'b1;
			partial_clause[7][114] 	= partial_clause_prev[7][114] & 1'b1;
			partial_clause[7][115] 	= partial_clause_prev[7][115] & 1'b1;
			partial_clause[7][116] 	= partial_clause_prev[7][116] & 1'b1;
			partial_clause[7][117] 	= partial_clause_prev[7][117] & 1'b1;
			partial_clause[7][118] 	= partial_clause_prev[7][118] & 1'b1;
			partial_clause[7][119] 	= partial_clause_prev[7][119] & 1'b1;
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & 1'b1;
			partial_clause[7][123] 	= partial_clause_prev[7][123] & 1'b1;
			partial_clause[7][124] 	= partial_clause_prev[7][124] & 1'b1;
			partial_clause[7][125] 	= partial_clause_prev[7][125] & 1'b1;
			partial_clause[7][126] 	= partial_clause_prev[7][126] & 1'b1;
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & 1'b1;
			partial_clause[7][129] 	= partial_clause_prev[7][129] & 1'b1;
			partial_clause[7][130] 	= partial_clause_prev[7][130] & 1'b1;
			partial_clause[7][131] 	= partial_clause_prev[7][131] & 1'b1;
			partial_clause[7][132] 	= partial_clause_prev[7][132] & 1'b1;
			partial_clause[7][133] 	= partial_clause_prev[7][133] & 1'b1;
			partial_clause[7][134] 	= partial_clause_prev[7][134] & 1'b1;
			partial_clause[7][135] 	= partial_clause_prev[7][135] & 1'b1;
			partial_clause[7][136] 	= partial_clause_prev[7][136] & 1'b1;
			partial_clause[7][137] 	= partial_clause_prev[7][137] & 1'b1;
			partial_clause[7][138] 	= partial_clause_prev[7][138] & 1'b1;
			partial_clause[7][139] 	= partial_clause_prev[7][139] & 1'b1;
			partial_clause[7][140] 	= partial_clause_prev[7][140] & 1'b1;
			partial_clause[7][141] 	= partial_clause_prev[7][141] & ~x[7];
			partial_clause[7][142] 	= partial_clause_prev[7][142] & 1'b1;
			partial_clause[7][143] 	= partial_clause_prev[7][143] & 1'b1;
			partial_clause[7][144] 	= partial_clause_prev[7][144] & 1'b1;
			partial_clause[7][145] 	= partial_clause_prev[7][145] & 1'b1;
			partial_clause[7][146] 	= partial_clause_prev[7][146] & 1'b1;
			partial_clause[7][147] 	= partial_clause_prev[7][147] & 1'b1;
			partial_clause[7][148] 	= partial_clause_prev[7][148] & 1'b1;
			partial_clause[7][149] 	= partial_clause_prev[7][149] & 1'b1;
			partial_clause[7][150] 	= partial_clause_prev[7][150] & 1'b1;
			partial_clause[7][151] 	= partial_clause_prev[7][151] & 1'b1;
			partial_clause[7][152] 	= partial_clause_prev[7][152] & 1'b1;
			partial_clause[7][153] 	= partial_clause_prev[7][153] & 1'b1;
			partial_clause[7][154] 	= partial_clause_prev[7][154] & 1'b1;
			partial_clause[7][155] 	= partial_clause_prev[7][155] & 1'b1;
			partial_clause[7][156] 	= partial_clause_prev[7][156] & 1'b1;
			partial_clause[7][157] 	= partial_clause_prev[7][157] & 1'b1;
			partial_clause[7][158] 	= partial_clause_prev[7][158] & 1'b1;
			partial_clause[7][159] 	= partial_clause_prev[7][159] & 1'b1;
			partial_clause[7][160] 	= partial_clause_prev[7][160] & 1'b1;
			partial_clause[7][161] 	= partial_clause_prev[7][161] & 1'b1;
			partial_clause[7][162] 	= partial_clause_prev[7][162] & 1'b1;
			partial_clause[7][163] 	= partial_clause_prev[7][163] & 1'b1;
			partial_clause[7][164] 	= partial_clause_prev[7][164] & 1'b1;
			partial_clause[7][165] 	= partial_clause_prev[7][165] & 1'b1;
			partial_clause[7][166] 	= partial_clause_prev[7][166] & ~x[44];
			partial_clause[7][167] 	= partial_clause_prev[7][167] & 1'b1;
			partial_clause[7][168] 	= partial_clause_prev[7][168] & 1'b1;
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & 1'b1;
			partial_clause[7][171] 	= partial_clause_prev[7][171] & 1'b1;
			partial_clause[7][172] 	= partial_clause_prev[7][172] & 1'b1;
			partial_clause[7][173] 	= partial_clause_prev[7][173] & 1'b1;
			partial_clause[7][174] 	= partial_clause_prev[7][174] & 1'b1;
			partial_clause[7][175] 	= partial_clause_prev[7][175] & 1'b1;
			partial_clause[7][176] 	= partial_clause_prev[7][176] & 1'b1;
			partial_clause[7][177] 	= partial_clause_prev[7][177] & 1'b1;
			partial_clause[7][178] 	= partial_clause_prev[7][178] & 1'b1;
			partial_clause[7][179] 	= partial_clause_prev[7][179] & 1'b1;
			partial_clause[7][180] 	= partial_clause_prev[7][180] & 1'b1;
			partial_clause[7][181] 	= partial_clause_prev[7][181] & 1'b1;
			partial_clause[7][182] 	= partial_clause_prev[7][182] & 1'b1;
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & 1'b1;
			partial_clause[7][185] 	= partial_clause_prev[7][185] & ~x[56];
			partial_clause[7][186] 	= partial_clause_prev[7][186] & 1'b1;
			partial_clause[7][187] 	= partial_clause_prev[7][187] & 1'b1;
			partial_clause[7][188] 	= partial_clause_prev[7][188] & 1'b1;
			partial_clause[7][189] 	= partial_clause_prev[7][189] & 1'b1;
			partial_clause[7][190] 	= partial_clause_prev[7][190] & 1'b1;
			partial_clause[7][191] 	= partial_clause_prev[7][191] & 1'b1;
			partial_clause[7][192] 	= partial_clause_prev[7][192] & 1'b1;
			partial_clause[7][193] 	= partial_clause_prev[7][193] & 1'b1;
			partial_clause[7][194] 	= partial_clause_prev[7][194] & 1'b1;
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & ~x[53];
			partial_clause[7][197] 	= partial_clause_prev[7][197] & 1'b1;
			partial_clause[7][198] 	= partial_clause_prev[7][198] & 1'b1;
			partial_clause[7][199] 	= partial_clause_prev[7][199] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & x[24];
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & x[32];
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & x[29];
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			partial_clause[8][100] 	= partial_clause_prev[8][100] & 1'b1;
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & 1'b1;
			partial_clause[8][103] 	= partial_clause_prev[8][103] & 1'b1;
			partial_clause[8][104] 	= partial_clause_prev[8][104] & 1'b1;
			partial_clause[8][105] 	= partial_clause_prev[8][105] & 1'b1;
			partial_clause[8][106] 	= partial_clause_prev[8][106] & 1'b1;
			partial_clause[8][107] 	= partial_clause_prev[8][107] & 1'b1;
			partial_clause[8][108] 	= partial_clause_prev[8][108] & 1'b1;
			partial_clause[8][109] 	= partial_clause_prev[8][109] & 1'b1;
			partial_clause[8][110] 	= partial_clause_prev[8][110] & 1'b1;
			partial_clause[8][111] 	= partial_clause_prev[8][111] & 1'b1;
			partial_clause[8][112] 	= partial_clause_prev[8][112] & 1'b1;
			partial_clause[8][113] 	= partial_clause_prev[8][113] & 1'b1;
			partial_clause[8][114] 	= partial_clause_prev[8][114] & 1'b1;
			partial_clause[8][115] 	= partial_clause_prev[8][115] & 1'b1;
			partial_clause[8][116] 	= partial_clause_prev[8][116] & 1'b1;
			partial_clause[8][117] 	= partial_clause_prev[8][117] & 1'b1;
			partial_clause[8][118] 	= partial_clause_prev[8][118] & 1'b1;
			partial_clause[8][119] 	= partial_clause_prev[8][119] & 1'b1;
			partial_clause[8][120] 	= partial_clause_prev[8][120] & 1'b1;
			partial_clause[8][121] 	= partial_clause_prev[8][121] & 1'b1;
			partial_clause[8][122] 	= partial_clause_prev[8][122] & 1'b1;
			partial_clause[8][123] 	= partial_clause_prev[8][123] & x[4];
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & 1'b1;
			partial_clause[8][126] 	= partial_clause_prev[8][126] & 1'b1;
			partial_clause[8][127] 	= partial_clause_prev[8][127] & 1'b1;
			partial_clause[8][128] 	= partial_clause_prev[8][128] & 1'b1;
			partial_clause[8][129] 	= partial_clause_prev[8][129] & 1'b1;
			partial_clause[8][130] 	= partial_clause_prev[8][130] & 1'b1;
			partial_clause[8][131] 	= partial_clause_prev[8][131] & 1'b1;
			partial_clause[8][132] 	= partial_clause_prev[8][132] & 1'b1;
			partial_clause[8][133] 	= partial_clause_prev[8][133] & 1'b1;
			partial_clause[8][134] 	= partial_clause_prev[8][134] & 1'b1;
			partial_clause[8][135] 	= partial_clause_prev[8][135] & ~x[9];
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & 1'b1;
			partial_clause[8][138] 	= partial_clause_prev[8][138] & 1'b1;
			partial_clause[8][139] 	= partial_clause_prev[8][139] & 1'b1;
			partial_clause[8][140] 	= partial_clause_prev[8][140] & 1'b1;
			partial_clause[8][141] 	= partial_clause_prev[8][141] & 1'b1;
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & 1'b1;
			partial_clause[8][144] 	= partial_clause_prev[8][144] & 1'b1;
			partial_clause[8][145] 	= partial_clause_prev[8][145] & 1'b1;
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & 1'b1;
			partial_clause[8][148] 	= partial_clause_prev[8][148] & 1'b1;
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & 1'b1;
			partial_clause[8][151] 	= partial_clause_prev[8][151] & 1'b1;
			partial_clause[8][152] 	= partial_clause_prev[8][152] & 1'b1;
			partial_clause[8][153] 	= partial_clause_prev[8][153] & 1'b1;
			partial_clause[8][154] 	= partial_clause_prev[8][154] & 1'b1;
			partial_clause[8][155] 	= partial_clause_prev[8][155] & 1'b1;
			partial_clause[8][156] 	= partial_clause_prev[8][156] & 1'b1;
			partial_clause[8][157] 	= partial_clause_prev[8][157] & x[22];
			partial_clause[8][158] 	= partial_clause_prev[8][158] & x[22];
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & 1'b1;
			partial_clause[8][161] 	= partial_clause_prev[8][161] & 1'b1;
			partial_clause[8][162] 	= partial_clause_prev[8][162] & 1'b1;
			partial_clause[8][163] 	= partial_clause_prev[8][163] & 1'b1;
			partial_clause[8][164] 	= partial_clause_prev[8][164] & 1'b1;
			partial_clause[8][165] 	= partial_clause_prev[8][165] & 1'b1;
			partial_clause[8][166] 	= partial_clause_prev[8][166] & 1'b1;
			partial_clause[8][167] 	= partial_clause_prev[8][167] & 1'b1;
			partial_clause[8][168] 	= partial_clause_prev[8][168] & 1'b1;
			partial_clause[8][169] 	= partial_clause_prev[8][169] & 1'b1;
			partial_clause[8][170] 	= partial_clause_prev[8][170] & 1'b1;
			partial_clause[8][171] 	= partial_clause_prev[8][171] & 1'b1;
			partial_clause[8][172] 	= partial_clause_prev[8][172] & 1'b1;
			partial_clause[8][173] 	= partial_clause_prev[8][173] & 1'b1;
			partial_clause[8][174] 	= partial_clause_prev[8][174] & x[37];
			partial_clause[8][175] 	= partial_clause_prev[8][175] & 1'b1;
			partial_clause[8][176] 	= partial_clause_prev[8][176] & 1'b1;
			partial_clause[8][177] 	= partial_clause_prev[8][177] & 1'b1;
			partial_clause[8][178] 	= partial_clause_prev[8][178] & 1'b1;
			partial_clause[8][179] 	= partial_clause_prev[8][179] & 1'b1;
			partial_clause[8][180] 	= partial_clause_prev[8][180] & 1'b1;
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & 1'b1;
			partial_clause[8][183] 	= partial_clause_prev[8][183] & 1'b1;
			partial_clause[8][184] 	= partial_clause_prev[8][184] & 1'b1;
			partial_clause[8][185] 	= partial_clause_prev[8][185] & 1'b1;
			partial_clause[8][186] 	= partial_clause_prev[8][186] & 1'b1;
			partial_clause[8][187] 	= partial_clause_prev[8][187] & 1'b1;
			partial_clause[8][188] 	= partial_clause_prev[8][188] & 1'b1;
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & 1'b1;
			partial_clause[8][191] 	= partial_clause_prev[8][191] & 1'b1;
			partial_clause[8][192] 	= partial_clause_prev[8][192] & 1'b1;
			partial_clause[8][193] 	= partial_clause_prev[8][193] & 1'b1;
			partial_clause[8][194] 	= partial_clause_prev[8][194] & 1'b1;
			partial_clause[8][195] 	= partial_clause_prev[8][195] & 1'b1;
			partial_clause[8][196] 	= partial_clause_prev[8][196] & 1'b1;
			partial_clause[8][197] 	= partial_clause_prev[8][197] & 1'b1;
			partial_clause[8][198] 	= partial_clause_prev[8][198] & x[7];
			partial_clause[8][199] 	= partial_clause_prev[8][199] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & x[15];
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & x[14];
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & x[15];
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & x[11];
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & x[17];
			partial_clause[9][20] 	= partial_clause_prev[9][20] & x[20];
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & x[14];
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & 1'b1;
			partial_clause[9][36] 	= partial_clause_prev[9][36] & x[18];
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & x[3];
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & x[18];
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & x[17];
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & x[14];
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & x[15];
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & x[16];
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & x[16];
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & x[13];
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
			partial_clause[9][100] 	= partial_clause_prev[9][100] & 1'b1;
			partial_clause[9][101] 	= partial_clause_prev[9][101] & ~x[13] & ~x[18];
			partial_clause[9][102] 	= partial_clause_prev[9][102] & 1'b1;
			partial_clause[9][103] 	= partial_clause_prev[9][103] & 1'b1;
			partial_clause[9][104] 	= partial_clause_prev[9][104] & 1'b1;
			partial_clause[9][105] 	= partial_clause_prev[9][105] & 1'b1;
			partial_clause[9][106] 	= partial_clause_prev[9][106] & 1'b1;
			partial_clause[9][107] 	= partial_clause_prev[9][107] & 1'b1;
			partial_clause[9][108] 	= partial_clause_prev[9][108] & 1'b1;
			partial_clause[9][109] 	= partial_clause_prev[9][109] & 1'b1;
			partial_clause[9][110] 	= partial_clause_prev[9][110] & 1'b1;
			partial_clause[9][111] 	= partial_clause_prev[9][111] & 1'b1;
			partial_clause[9][112] 	= partial_clause_prev[9][112] & 1'b1;
			partial_clause[9][113] 	= partial_clause_prev[9][113] & 1'b1;
			partial_clause[9][114] 	= partial_clause_prev[9][114] & 1'b1;
			partial_clause[9][115] 	= partial_clause_prev[9][115] & 1'b1;
			partial_clause[9][116] 	= partial_clause_prev[9][116] & 1'b1;
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & 1'b1;
			partial_clause[9][119] 	= partial_clause_prev[9][119] & 1'b1;
			partial_clause[9][120] 	= partial_clause_prev[9][120] & 1'b1;
			partial_clause[9][121] 	= partial_clause_prev[9][121] & 1'b1;
			partial_clause[9][122] 	= partial_clause_prev[9][122] & 1'b1;
			partial_clause[9][123] 	= partial_clause_prev[9][123] & 1'b1;
			partial_clause[9][124] 	= partial_clause_prev[9][124] & 1'b1;
			partial_clause[9][125] 	= partial_clause_prev[9][125] & 1'b1;
			partial_clause[9][126] 	= partial_clause_prev[9][126] & 1'b1;
			partial_clause[9][127] 	= partial_clause_prev[9][127] & 1'b1;
			partial_clause[9][128] 	= partial_clause_prev[9][128] & 1'b1;
			partial_clause[9][129] 	= partial_clause_prev[9][129] & 1'b1;
			partial_clause[9][130] 	= partial_clause_prev[9][130] & 1'b1;
			partial_clause[9][131] 	= partial_clause_prev[9][131] & 1'b1;
			partial_clause[9][132] 	= partial_clause_prev[9][132] & 1'b1;
			partial_clause[9][133] 	= partial_clause_prev[9][133] & 1'b1;
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & 1'b1;
			partial_clause[9][138] 	= partial_clause_prev[9][138] & 1'b1;
			partial_clause[9][139] 	= partial_clause_prev[9][139] & 1'b1;
			partial_clause[9][140] 	= partial_clause_prev[9][140] & 1'b1;
			partial_clause[9][141] 	= partial_clause_prev[9][141] & 1'b1;
			partial_clause[9][142] 	= partial_clause_prev[9][142] & 1'b1;
			partial_clause[9][143] 	= partial_clause_prev[9][143] & 1'b1;
			partial_clause[9][144] 	= partial_clause_prev[9][144] & 1'b1;
			partial_clause[9][145] 	= partial_clause_prev[9][145] & 1'b1;
			partial_clause[9][146] 	= partial_clause_prev[9][146] & 1'b1;
			partial_clause[9][147] 	= partial_clause_prev[9][147] & 1'b1;
			partial_clause[9][148] 	= partial_clause_prev[9][148] & 1'b1;
			partial_clause[9][149] 	= partial_clause_prev[9][149] & 1'b1;
			partial_clause[9][150] 	= partial_clause_prev[9][150] & 1'b1;
			partial_clause[9][151] 	= partial_clause_prev[9][151] & ~x[8];
			partial_clause[9][152] 	= partial_clause_prev[9][152] & 1'b1;
			partial_clause[9][153] 	= partial_clause_prev[9][153] & 1'b1;
			partial_clause[9][154] 	= partial_clause_prev[9][154] & 1'b1;
			partial_clause[9][155] 	= partial_clause_prev[9][155] & 1'b1;
			partial_clause[9][156] 	= partial_clause_prev[9][156] & 1'b1;
			partial_clause[9][157] 	= partial_clause_prev[9][157] & 1'b1;
			partial_clause[9][158] 	= partial_clause_prev[9][158] & 1'b1;
			partial_clause[9][159] 	= partial_clause_prev[9][159] & 1'b1;
			partial_clause[9][160] 	= partial_clause_prev[9][160] & 1'b1;
			partial_clause[9][161] 	= partial_clause_prev[9][161] & 1'b1;
			partial_clause[9][162] 	= partial_clause_prev[9][162] & 1'b1;
			partial_clause[9][163] 	= partial_clause_prev[9][163] & 1'b1;
			partial_clause[9][164] 	= partial_clause_prev[9][164] & 1'b1;
			partial_clause[9][165] 	= partial_clause_prev[9][165] & 1'b1;
			partial_clause[9][166] 	= partial_clause_prev[9][166] & 1'b1;
			partial_clause[9][167] 	= partial_clause_prev[9][167] & 1'b1;
			partial_clause[9][168] 	= partial_clause_prev[9][168] & ~x[7];
			partial_clause[9][169] 	= partial_clause_prev[9][169] & 1'b1;
			partial_clause[9][170] 	= partial_clause_prev[9][170] & 1'b1;
			partial_clause[9][171] 	= partial_clause_prev[9][171] & 1'b1;
			partial_clause[9][172] 	= partial_clause_prev[9][172] & 1'b1;
			partial_clause[9][173] 	= partial_clause_prev[9][173] & 1'b1;
			partial_clause[9][174] 	= partial_clause_prev[9][174] & 1'b1;
			partial_clause[9][175] 	= partial_clause_prev[9][175] & 1'b1;
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & 1'b1;
			partial_clause[9][178] 	= partial_clause_prev[9][178] & 1'b1;
			partial_clause[9][179] 	= partial_clause_prev[9][179] & 1'b1;
			partial_clause[9][180] 	= partial_clause_prev[9][180] & 1'b1;
			partial_clause[9][181] 	= partial_clause_prev[9][181] & 1'b1;
			partial_clause[9][182] 	= partial_clause_prev[9][182] & 1'b1;
			partial_clause[9][183] 	= partial_clause_prev[9][183] & 1'b1;
			partial_clause[9][184] 	= partial_clause_prev[9][184] & 1'b1;
			partial_clause[9][185] 	= partial_clause_prev[9][185] & 1'b1;
			partial_clause[9][186] 	= partial_clause_prev[9][186] & 1'b1;
			partial_clause[9][187] 	= partial_clause_prev[9][187] & 1'b1;
			partial_clause[9][188] 	= partial_clause_prev[9][188] & 1'b1;
			partial_clause[9][189] 	= partial_clause_prev[9][189] & 1'b1;
			partial_clause[9][190] 	= partial_clause_prev[9][190] & 1'b1;
			partial_clause[9][191] 	= partial_clause_prev[9][191] & 1'b1;
			partial_clause[9][192] 	= partial_clause_prev[9][192] & 1'b1;
			partial_clause[9][193] 	= partial_clause_prev[9][193] & 1'b1;
			partial_clause[9][194] 	= partial_clause_prev[9][194] & 1'b1;
			partial_clause[9][195] 	= partial_clause_prev[9][195] & 1'b1;
			partial_clause[9][196] 	= partial_clause_prev[9][196] & 1'b1;
			partial_clause[9][197] 	= partial_clause_prev[9][197] & 1'b1;
			partial_clause[9][198] 	= partial_clause_prev[9][198] & 1'b1;
			partial_clause[9][199] 	= partial_clause_prev[9][199] & 1'b1;
		end
	end
endmodule


module HCB_12 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [199:0] partial_clause_prev [10];
	output	logic[199:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & x[6];
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & x[2];
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			partial_clause[0][100] 	= partial_clause_prev[0][100] & 1'b1;
			partial_clause[0][101] 	= partial_clause_prev[0][101] & 1'b1;
			partial_clause[0][102] 	= partial_clause_prev[0][102] & 1'b1;
			partial_clause[0][103] 	= partial_clause_prev[0][103] & 1'b1;
			partial_clause[0][104] 	= partial_clause_prev[0][104] & 1'b1;
			partial_clause[0][105] 	= partial_clause_prev[0][105] & 1'b1;
			partial_clause[0][106] 	= partial_clause_prev[0][106] & 1'b1;
			partial_clause[0][107] 	= partial_clause_prev[0][107] & 1'b1;
			partial_clause[0][108] 	= partial_clause_prev[0][108] & 1'b1;
			partial_clause[0][109] 	= partial_clause_prev[0][109] & 1'b1;
			partial_clause[0][110] 	= partial_clause_prev[0][110] & 1'b1;
			partial_clause[0][111] 	= partial_clause_prev[0][111] & 1'b1;
			partial_clause[0][112] 	= partial_clause_prev[0][112] & 1'b1;
			partial_clause[0][113] 	= partial_clause_prev[0][113] & 1'b1;
			partial_clause[0][114] 	= partial_clause_prev[0][114] & 1'b1;
			partial_clause[0][115] 	= partial_clause_prev[0][115] & 1'b1;
			partial_clause[0][116] 	= partial_clause_prev[0][116] & 1'b1;
			partial_clause[0][117] 	= partial_clause_prev[0][117] & 1'b1;
			partial_clause[0][118] 	= partial_clause_prev[0][118] & 1'b1;
			partial_clause[0][119] 	= partial_clause_prev[0][119] & 1'b1;
			partial_clause[0][120] 	= partial_clause_prev[0][120] & 1'b1;
			partial_clause[0][121] 	= partial_clause_prev[0][121] & 1'b1;
			partial_clause[0][122] 	= partial_clause_prev[0][122] & 1'b1;
			partial_clause[0][123] 	= partial_clause_prev[0][123] & 1'b1;
			partial_clause[0][124] 	= partial_clause_prev[0][124] & 1'b1;
			partial_clause[0][125] 	= partial_clause_prev[0][125] & 1'b1;
			partial_clause[0][126] 	= partial_clause_prev[0][126] & 1'b1;
			partial_clause[0][127] 	= partial_clause_prev[0][127] & 1'b1;
			partial_clause[0][128] 	= partial_clause_prev[0][128] & 1'b1;
			partial_clause[0][129] 	= partial_clause_prev[0][129] & 1'b1;
			partial_clause[0][130] 	= partial_clause_prev[0][130] & 1'b1;
			partial_clause[0][131] 	= partial_clause_prev[0][131] & 1'b1;
			partial_clause[0][132] 	= partial_clause_prev[0][132] & 1'b1;
			partial_clause[0][133] 	= partial_clause_prev[0][133] & 1'b1;
			partial_clause[0][134] 	= partial_clause_prev[0][134] & 1'b1;
			partial_clause[0][135] 	= partial_clause_prev[0][135] & 1'b1;
			partial_clause[0][136] 	= partial_clause_prev[0][136] & 1'b1;
			partial_clause[0][137] 	= partial_clause_prev[0][137] & 1'b1;
			partial_clause[0][138] 	= partial_clause_prev[0][138] & 1'b1;
			partial_clause[0][139] 	= partial_clause_prev[0][139] & 1'b1;
			partial_clause[0][140] 	= partial_clause_prev[0][140] & 1'b1;
			partial_clause[0][141] 	= partial_clause_prev[0][141] & 1'b1;
			partial_clause[0][142] 	= partial_clause_prev[0][142] & 1'b1;
			partial_clause[0][143] 	= partial_clause_prev[0][143] & 1'b1;
			partial_clause[0][144] 	= partial_clause_prev[0][144] & 1'b1;
			partial_clause[0][145] 	= partial_clause_prev[0][145] & 1'b1;
			partial_clause[0][146] 	= partial_clause_prev[0][146] & 1'b1;
			partial_clause[0][147] 	= partial_clause_prev[0][147] & 1'b1;
			partial_clause[0][148] 	= partial_clause_prev[0][148] & 1'b1;
			partial_clause[0][149] 	= partial_clause_prev[0][149] & 1'b1;
			partial_clause[0][150] 	= partial_clause_prev[0][150] & 1'b1;
			partial_clause[0][151] 	= partial_clause_prev[0][151] & 1'b1;
			partial_clause[0][152] 	= partial_clause_prev[0][152] & 1'b1;
			partial_clause[0][153] 	= partial_clause_prev[0][153] & 1'b1;
			partial_clause[0][154] 	= partial_clause_prev[0][154] & 1'b1;
			partial_clause[0][155] 	= partial_clause_prev[0][155] & 1'b1;
			partial_clause[0][156] 	= partial_clause_prev[0][156] & 1'b1;
			partial_clause[0][157] 	= partial_clause_prev[0][157] & 1'b1;
			partial_clause[0][158] 	= partial_clause_prev[0][158] & 1'b1;
			partial_clause[0][159] 	= partial_clause_prev[0][159] & 1'b1;
			partial_clause[0][160] 	= partial_clause_prev[0][160] & 1'b1;
			partial_clause[0][161] 	= partial_clause_prev[0][161] & 1'b1;
			partial_clause[0][162] 	= partial_clause_prev[0][162] & 1'b1;
			partial_clause[0][163] 	= partial_clause_prev[0][163] & 1'b1;
			partial_clause[0][164] 	= partial_clause_prev[0][164] & 1'b1;
			partial_clause[0][165] 	= partial_clause_prev[0][165] & 1'b1;
			partial_clause[0][166] 	= partial_clause_prev[0][166] & 1'b1;
			partial_clause[0][167] 	= partial_clause_prev[0][167] & 1'b1;
			partial_clause[0][168] 	= partial_clause_prev[0][168] & 1'b1;
			partial_clause[0][169] 	= partial_clause_prev[0][169] & 1'b1;
			partial_clause[0][170] 	= partial_clause_prev[0][170] & 1'b1;
			partial_clause[0][171] 	= partial_clause_prev[0][171] & 1'b1;
			partial_clause[0][172] 	= partial_clause_prev[0][172] & 1'b1;
			partial_clause[0][173] 	= partial_clause_prev[0][173] & 1'b1;
			partial_clause[0][174] 	= partial_clause_prev[0][174] & 1'b1;
			partial_clause[0][175] 	= partial_clause_prev[0][175] & 1'b1;
			partial_clause[0][176] 	= partial_clause_prev[0][176] & 1'b1;
			partial_clause[0][177] 	= partial_clause_prev[0][177] & 1'b1;
			partial_clause[0][178] 	= partial_clause_prev[0][178] & 1'b1;
			partial_clause[0][179] 	= partial_clause_prev[0][179] & 1'b1;
			partial_clause[0][180] 	= partial_clause_prev[0][180] & 1'b1;
			partial_clause[0][181] 	= partial_clause_prev[0][181] & 1'b1;
			partial_clause[0][182] 	= partial_clause_prev[0][182] & 1'b1;
			partial_clause[0][183] 	= partial_clause_prev[0][183] & 1'b1;
			partial_clause[0][184] 	= partial_clause_prev[0][184] & 1'b1;
			partial_clause[0][185] 	= partial_clause_prev[0][185] & 1'b1;
			partial_clause[0][186] 	= partial_clause_prev[0][186] & 1'b1;
			partial_clause[0][187] 	= partial_clause_prev[0][187] & 1'b1;
			partial_clause[0][188] 	= partial_clause_prev[0][188] & 1'b1;
			partial_clause[0][189] 	= partial_clause_prev[0][189] & 1'b1;
			partial_clause[0][190] 	= partial_clause_prev[0][190] & 1'b1;
			partial_clause[0][191] 	= partial_clause_prev[0][191] & 1'b1;
			partial_clause[0][192] 	= partial_clause_prev[0][192] & 1'b1;
			partial_clause[0][193] 	= partial_clause_prev[0][193] & 1'b1;
			partial_clause[0][194] 	= partial_clause_prev[0][194] & 1'b1;
			partial_clause[0][195] 	= partial_clause_prev[0][195] & 1'b1;
			partial_clause[0][196] 	= partial_clause_prev[0][196] & 1'b1;
			partial_clause[0][197] 	= partial_clause_prev[0][197] & 1'b1;
			partial_clause[0][198] 	= partial_clause_prev[0][198] & 1'b1;
			partial_clause[0][199] 	= partial_clause_prev[0][199] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & x[11];
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & x[7];
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & 1'b1;
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & 1'b1;
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & x[9];
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			partial_clause[1][100] 	= partial_clause_prev[1][100] & 1'b1;
			partial_clause[1][101] 	= partial_clause_prev[1][101] & 1'b1;
			partial_clause[1][102] 	= partial_clause_prev[1][102] & 1'b1;
			partial_clause[1][103] 	= partial_clause_prev[1][103] & 1'b1;
			partial_clause[1][104] 	= partial_clause_prev[1][104] & 1'b1;
			partial_clause[1][105] 	= partial_clause_prev[1][105] & 1'b1;
			partial_clause[1][106] 	= partial_clause_prev[1][106] & 1'b1;
			partial_clause[1][107] 	= partial_clause_prev[1][107] & 1'b1;
			partial_clause[1][108] 	= partial_clause_prev[1][108] & 1'b1;
			partial_clause[1][109] 	= partial_clause_prev[1][109] & 1'b1;
			partial_clause[1][110] 	= partial_clause_prev[1][110] & 1'b1;
			partial_clause[1][111] 	= partial_clause_prev[1][111] & 1'b1;
			partial_clause[1][112] 	= partial_clause_prev[1][112] & 1'b1;
			partial_clause[1][113] 	= partial_clause_prev[1][113] & 1'b1;
			partial_clause[1][114] 	= partial_clause_prev[1][114] & 1'b1;
			partial_clause[1][115] 	= partial_clause_prev[1][115] & 1'b1;
			partial_clause[1][116] 	= partial_clause_prev[1][116] & 1'b1;
			partial_clause[1][117] 	= partial_clause_prev[1][117] & 1'b1;
			partial_clause[1][118] 	= partial_clause_prev[1][118] & 1'b1;
			partial_clause[1][119] 	= partial_clause_prev[1][119] & 1'b1;
			partial_clause[1][120] 	= partial_clause_prev[1][120] & 1'b1;
			partial_clause[1][121] 	= partial_clause_prev[1][121] & 1'b1;
			partial_clause[1][122] 	= partial_clause_prev[1][122] & 1'b1;
			partial_clause[1][123] 	= partial_clause_prev[1][123] & 1'b1;
			partial_clause[1][124] 	= partial_clause_prev[1][124] & 1'b1;
			partial_clause[1][125] 	= partial_clause_prev[1][125] & 1'b1;
			partial_clause[1][126] 	= partial_clause_prev[1][126] & 1'b1;
			partial_clause[1][127] 	= partial_clause_prev[1][127] & 1'b1;
			partial_clause[1][128] 	= partial_clause_prev[1][128] & 1'b1;
			partial_clause[1][129] 	= partial_clause_prev[1][129] & 1'b1;
			partial_clause[1][130] 	= partial_clause_prev[1][130] & 1'b1;
			partial_clause[1][131] 	= partial_clause_prev[1][131] & 1'b1;
			partial_clause[1][132] 	= partial_clause_prev[1][132] & 1'b1;
			partial_clause[1][133] 	= partial_clause_prev[1][133] & 1'b1;
			partial_clause[1][134] 	= partial_clause_prev[1][134] & 1'b1;
			partial_clause[1][135] 	= partial_clause_prev[1][135] & 1'b1;
			partial_clause[1][136] 	= partial_clause_prev[1][136] & 1'b1;
			partial_clause[1][137] 	= partial_clause_prev[1][137] & 1'b1;
			partial_clause[1][138] 	= partial_clause_prev[1][138] & 1'b1;
			partial_clause[1][139] 	= partial_clause_prev[1][139] & 1'b1;
			partial_clause[1][140] 	= partial_clause_prev[1][140] & 1'b1;
			partial_clause[1][141] 	= partial_clause_prev[1][141] & 1'b1;
			partial_clause[1][142] 	= partial_clause_prev[1][142] & 1'b1;
			partial_clause[1][143] 	= partial_clause_prev[1][143] & 1'b1;
			partial_clause[1][144] 	= partial_clause_prev[1][144] & 1'b1;
			partial_clause[1][145] 	= partial_clause_prev[1][145] & 1'b1;
			partial_clause[1][146] 	= partial_clause_prev[1][146] & 1'b1;
			partial_clause[1][147] 	= partial_clause_prev[1][147] & 1'b1;
			partial_clause[1][148] 	= partial_clause_prev[1][148] & 1'b1;
			partial_clause[1][149] 	= partial_clause_prev[1][149] & 1'b1;
			partial_clause[1][150] 	= partial_clause_prev[1][150] & 1'b1;
			partial_clause[1][151] 	= partial_clause_prev[1][151] & 1'b1;
			partial_clause[1][152] 	= partial_clause_prev[1][152] & 1'b1;
			partial_clause[1][153] 	= partial_clause_prev[1][153] & 1'b1;
			partial_clause[1][154] 	= partial_clause_prev[1][154] & 1'b1;
			partial_clause[1][155] 	= partial_clause_prev[1][155] & 1'b1;
			partial_clause[1][156] 	= partial_clause_prev[1][156] & 1'b1;
			partial_clause[1][157] 	= partial_clause_prev[1][157] & 1'b1;
			partial_clause[1][158] 	= partial_clause_prev[1][158] & 1'b1;
			partial_clause[1][159] 	= partial_clause_prev[1][159] & 1'b1;
			partial_clause[1][160] 	= partial_clause_prev[1][160] & 1'b1;
			partial_clause[1][161] 	= partial_clause_prev[1][161] & 1'b1;
			partial_clause[1][162] 	= partial_clause_prev[1][162] & 1'b1;
			partial_clause[1][163] 	= partial_clause_prev[1][163] & 1'b1;
			partial_clause[1][164] 	= partial_clause_prev[1][164] & 1'b1;
			partial_clause[1][165] 	= partial_clause_prev[1][165] & 1'b1;
			partial_clause[1][166] 	= partial_clause_prev[1][166] & 1'b1;
			partial_clause[1][167] 	= partial_clause_prev[1][167] & 1'b1;
			partial_clause[1][168] 	= partial_clause_prev[1][168] & 1'b1;
			partial_clause[1][169] 	= partial_clause_prev[1][169] & 1'b1;
			partial_clause[1][170] 	= partial_clause_prev[1][170] & 1'b1;
			partial_clause[1][171] 	= partial_clause_prev[1][171] & 1'b1;
			partial_clause[1][172] 	= partial_clause_prev[1][172] & 1'b1;
			partial_clause[1][173] 	= partial_clause_prev[1][173] & 1'b1;
			partial_clause[1][174] 	= partial_clause_prev[1][174] & 1'b1;
			partial_clause[1][175] 	= partial_clause_prev[1][175] & 1'b1;
			partial_clause[1][176] 	= partial_clause_prev[1][176] & 1'b1;
			partial_clause[1][177] 	= partial_clause_prev[1][177] & 1'b1;
			partial_clause[1][178] 	= partial_clause_prev[1][178] & 1'b1;
			partial_clause[1][179] 	= partial_clause_prev[1][179] & 1'b1;
			partial_clause[1][180] 	= partial_clause_prev[1][180] & 1'b1;
			partial_clause[1][181] 	= partial_clause_prev[1][181] & 1'b1;
			partial_clause[1][182] 	= partial_clause_prev[1][182] & 1'b1;
			partial_clause[1][183] 	= partial_clause_prev[1][183] & 1'b1;
			partial_clause[1][184] 	= partial_clause_prev[1][184] & 1'b1;
			partial_clause[1][185] 	= partial_clause_prev[1][185] & 1'b1;
			partial_clause[1][186] 	= partial_clause_prev[1][186] & 1'b1;
			partial_clause[1][187] 	= partial_clause_prev[1][187] & 1'b1;
			partial_clause[1][188] 	= partial_clause_prev[1][188] & 1'b1;
			partial_clause[1][189] 	= partial_clause_prev[1][189] & 1'b1;
			partial_clause[1][190] 	= partial_clause_prev[1][190] & 1'b1;
			partial_clause[1][191] 	= partial_clause_prev[1][191] & 1'b1;
			partial_clause[1][192] 	= partial_clause_prev[1][192] & 1'b1;
			partial_clause[1][193] 	= partial_clause_prev[1][193] & 1'b1;
			partial_clause[1][194] 	= partial_clause_prev[1][194] & 1'b1;
			partial_clause[1][195] 	= partial_clause_prev[1][195] & 1'b1;
			partial_clause[1][196] 	= partial_clause_prev[1][196] & 1'b1;
			partial_clause[1][197] 	= partial_clause_prev[1][197] & 1'b1;
			partial_clause[1][198] 	= partial_clause_prev[1][198] & 1'b1;
			partial_clause[1][199] 	= partial_clause_prev[1][199] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & 1'b1;
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			partial_clause[2][100] 	= partial_clause_prev[2][100] & 1'b1;
			partial_clause[2][101] 	= partial_clause_prev[2][101] & 1'b1;
			partial_clause[2][102] 	= partial_clause_prev[2][102] & 1'b1;
			partial_clause[2][103] 	= partial_clause_prev[2][103] & 1'b1;
			partial_clause[2][104] 	= partial_clause_prev[2][104] & 1'b1;
			partial_clause[2][105] 	= partial_clause_prev[2][105] & 1'b1;
			partial_clause[2][106] 	= partial_clause_prev[2][106] & 1'b1;
			partial_clause[2][107] 	= partial_clause_prev[2][107] & 1'b1;
			partial_clause[2][108] 	= partial_clause_prev[2][108] & 1'b1;
			partial_clause[2][109] 	= partial_clause_prev[2][109] & 1'b1;
			partial_clause[2][110] 	= partial_clause_prev[2][110] & 1'b1;
			partial_clause[2][111] 	= partial_clause_prev[2][111] & 1'b1;
			partial_clause[2][112] 	= partial_clause_prev[2][112] & 1'b1;
			partial_clause[2][113] 	= partial_clause_prev[2][113] & 1'b1;
			partial_clause[2][114] 	= partial_clause_prev[2][114] & 1'b1;
			partial_clause[2][115] 	= partial_clause_prev[2][115] & 1'b1;
			partial_clause[2][116] 	= partial_clause_prev[2][116] & 1'b1;
			partial_clause[2][117] 	= partial_clause_prev[2][117] & 1'b1;
			partial_clause[2][118] 	= partial_clause_prev[2][118] & 1'b1;
			partial_clause[2][119] 	= partial_clause_prev[2][119] & 1'b1;
			partial_clause[2][120] 	= partial_clause_prev[2][120] & 1'b1;
			partial_clause[2][121] 	= partial_clause_prev[2][121] & 1'b1;
			partial_clause[2][122] 	= partial_clause_prev[2][122] & 1'b1;
			partial_clause[2][123] 	= partial_clause_prev[2][123] & 1'b1;
			partial_clause[2][124] 	= partial_clause_prev[2][124] & 1'b1;
			partial_clause[2][125] 	= partial_clause_prev[2][125] & 1'b1;
			partial_clause[2][126] 	= partial_clause_prev[2][126] & 1'b1;
			partial_clause[2][127] 	= partial_clause_prev[2][127] & 1'b1;
			partial_clause[2][128] 	= partial_clause_prev[2][128] & 1'b1;
			partial_clause[2][129] 	= partial_clause_prev[2][129] & 1'b1;
			partial_clause[2][130] 	= partial_clause_prev[2][130] & 1'b1;
			partial_clause[2][131] 	= partial_clause_prev[2][131] & 1'b1;
			partial_clause[2][132] 	= partial_clause_prev[2][132] & 1'b1;
			partial_clause[2][133] 	= partial_clause_prev[2][133] & 1'b1;
			partial_clause[2][134] 	= partial_clause_prev[2][134] & 1'b1;
			partial_clause[2][135] 	= partial_clause_prev[2][135] & 1'b1;
			partial_clause[2][136] 	= partial_clause_prev[2][136] & 1'b1;
			partial_clause[2][137] 	= partial_clause_prev[2][137] & 1'b1;
			partial_clause[2][138] 	= partial_clause_prev[2][138] & 1'b1;
			partial_clause[2][139] 	= partial_clause_prev[2][139] & 1'b1;
			partial_clause[2][140] 	= partial_clause_prev[2][140] & 1'b1;
			partial_clause[2][141] 	= partial_clause_prev[2][141] & 1'b1;
			partial_clause[2][142] 	= partial_clause_prev[2][142] & 1'b1;
			partial_clause[2][143] 	= partial_clause_prev[2][143] & 1'b1;
			partial_clause[2][144] 	= partial_clause_prev[2][144] & 1'b1;
			partial_clause[2][145] 	= partial_clause_prev[2][145] & 1'b1;
			partial_clause[2][146] 	= partial_clause_prev[2][146] & 1'b1;
			partial_clause[2][147] 	= partial_clause_prev[2][147] & 1'b1;
			partial_clause[2][148] 	= partial_clause_prev[2][148] & 1'b1;
			partial_clause[2][149] 	= partial_clause_prev[2][149] & 1'b1;
			partial_clause[2][150] 	= partial_clause_prev[2][150] & 1'b1;
			partial_clause[2][151] 	= partial_clause_prev[2][151] & 1'b1;
			partial_clause[2][152] 	= partial_clause_prev[2][152] & 1'b1;
			partial_clause[2][153] 	= partial_clause_prev[2][153] & 1'b1;
			partial_clause[2][154] 	= partial_clause_prev[2][154] & 1'b1;
			partial_clause[2][155] 	= partial_clause_prev[2][155] & 1'b1;
			partial_clause[2][156] 	= partial_clause_prev[2][156] & 1'b1;
			partial_clause[2][157] 	= partial_clause_prev[2][157] & 1'b1;
			partial_clause[2][158] 	= partial_clause_prev[2][158] & 1'b1;
			partial_clause[2][159] 	= partial_clause_prev[2][159] & 1'b1;
			partial_clause[2][160] 	= partial_clause_prev[2][160] & 1'b1;
			partial_clause[2][161] 	= partial_clause_prev[2][161] & 1'b1;
			partial_clause[2][162] 	= partial_clause_prev[2][162] & 1'b1;
			partial_clause[2][163] 	= partial_clause_prev[2][163] & 1'b1;
			partial_clause[2][164] 	= partial_clause_prev[2][164] & 1'b1;
			partial_clause[2][165] 	= partial_clause_prev[2][165] & 1'b1;
			partial_clause[2][166] 	= partial_clause_prev[2][166] & 1'b1;
			partial_clause[2][167] 	= partial_clause_prev[2][167] & 1'b1;
			partial_clause[2][168] 	= partial_clause_prev[2][168] & 1'b1;
			partial_clause[2][169] 	= partial_clause_prev[2][169] & 1'b1;
			partial_clause[2][170] 	= partial_clause_prev[2][170] & 1'b1;
			partial_clause[2][171] 	= partial_clause_prev[2][171] & 1'b1;
			partial_clause[2][172] 	= partial_clause_prev[2][172] & 1'b1;
			partial_clause[2][173] 	= partial_clause_prev[2][173] & 1'b1;
			partial_clause[2][174] 	= partial_clause_prev[2][174] & 1'b1;
			partial_clause[2][175] 	= partial_clause_prev[2][175] & 1'b1;
			partial_clause[2][176] 	= partial_clause_prev[2][176] & 1'b1;
			partial_clause[2][177] 	= partial_clause_prev[2][177] & 1'b1;
			partial_clause[2][178] 	= partial_clause_prev[2][178] & 1'b1;
			partial_clause[2][179] 	= partial_clause_prev[2][179] & 1'b1;
			partial_clause[2][180] 	= partial_clause_prev[2][180] & 1'b1;
			partial_clause[2][181] 	= partial_clause_prev[2][181] & 1'b1;
			partial_clause[2][182] 	= partial_clause_prev[2][182] & 1'b1;
			partial_clause[2][183] 	= partial_clause_prev[2][183] & 1'b1;
			partial_clause[2][184] 	= partial_clause_prev[2][184] & 1'b1;
			partial_clause[2][185] 	= partial_clause_prev[2][185] & 1'b1;
			partial_clause[2][186] 	= partial_clause_prev[2][186] & 1'b1;
			partial_clause[2][187] 	= partial_clause_prev[2][187] & 1'b1;
			partial_clause[2][188] 	= partial_clause_prev[2][188] & 1'b1;
			partial_clause[2][189] 	= partial_clause_prev[2][189] & 1'b1;
			partial_clause[2][190] 	= partial_clause_prev[2][190] & 1'b1;
			partial_clause[2][191] 	= partial_clause_prev[2][191] & 1'b1;
			partial_clause[2][192] 	= partial_clause_prev[2][192] & 1'b1;
			partial_clause[2][193] 	= partial_clause_prev[2][193] & 1'b1;
			partial_clause[2][194] 	= partial_clause_prev[2][194] & 1'b1;
			partial_clause[2][195] 	= partial_clause_prev[2][195] & 1'b1;
			partial_clause[2][196] 	= partial_clause_prev[2][196] & 1'b1;
			partial_clause[2][197] 	= partial_clause_prev[2][197] & 1'b1;
			partial_clause[2][198] 	= partial_clause_prev[2][198] & 1'b1;
			partial_clause[2][199] 	= partial_clause_prev[2][199] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & x[4];
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & x[14];
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & x[14];
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & x[12];
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & 1'b1;
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			partial_clause[3][100] 	= partial_clause_prev[3][100] & 1'b1;
			partial_clause[3][101] 	= partial_clause_prev[3][101] & 1'b1;
			partial_clause[3][102] 	= partial_clause_prev[3][102] & 1'b1;
			partial_clause[3][103] 	= partial_clause_prev[3][103] & 1'b1;
			partial_clause[3][104] 	= partial_clause_prev[3][104] & 1'b1;
			partial_clause[3][105] 	= partial_clause_prev[3][105] & 1'b1;
			partial_clause[3][106] 	= partial_clause_prev[3][106] & 1'b1;
			partial_clause[3][107] 	= partial_clause_prev[3][107] & 1'b1;
			partial_clause[3][108] 	= partial_clause_prev[3][108] & 1'b1;
			partial_clause[3][109] 	= partial_clause_prev[3][109] & 1'b1;
			partial_clause[3][110] 	= partial_clause_prev[3][110] & 1'b1;
			partial_clause[3][111] 	= partial_clause_prev[3][111] & 1'b1;
			partial_clause[3][112] 	= partial_clause_prev[3][112] & 1'b1;
			partial_clause[3][113] 	= partial_clause_prev[3][113] & 1'b1;
			partial_clause[3][114] 	= partial_clause_prev[3][114] & 1'b1;
			partial_clause[3][115] 	= partial_clause_prev[3][115] & 1'b1;
			partial_clause[3][116] 	= partial_clause_prev[3][116] & 1'b1;
			partial_clause[3][117] 	= partial_clause_prev[3][117] & 1'b1;
			partial_clause[3][118] 	= partial_clause_prev[3][118] & 1'b1;
			partial_clause[3][119] 	= partial_clause_prev[3][119] & 1'b1;
			partial_clause[3][120] 	= partial_clause_prev[3][120] & 1'b1;
			partial_clause[3][121] 	= partial_clause_prev[3][121] & 1'b1;
			partial_clause[3][122] 	= partial_clause_prev[3][122] & 1'b1;
			partial_clause[3][123] 	= partial_clause_prev[3][123] & 1'b1;
			partial_clause[3][124] 	= partial_clause_prev[3][124] & 1'b1;
			partial_clause[3][125] 	= partial_clause_prev[3][125] & 1'b1;
			partial_clause[3][126] 	= partial_clause_prev[3][126] & 1'b1;
			partial_clause[3][127] 	= partial_clause_prev[3][127] & 1'b1;
			partial_clause[3][128] 	= partial_clause_prev[3][128] & 1'b1;
			partial_clause[3][129] 	= partial_clause_prev[3][129] & 1'b1;
			partial_clause[3][130] 	= partial_clause_prev[3][130] & 1'b1;
			partial_clause[3][131] 	= partial_clause_prev[3][131] & 1'b1;
			partial_clause[3][132] 	= partial_clause_prev[3][132] & 1'b1;
			partial_clause[3][133] 	= partial_clause_prev[3][133] & 1'b1;
			partial_clause[3][134] 	= partial_clause_prev[3][134] & 1'b1;
			partial_clause[3][135] 	= partial_clause_prev[3][135] & 1'b1;
			partial_clause[3][136] 	= partial_clause_prev[3][136] & 1'b1;
			partial_clause[3][137] 	= partial_clause_prev[3][137] & 1'b1;
			partial_clause[3][138] 	= partial_clause_prev[3][138] & 1'b1;
			partial_clause[3][139] 	= partial_clause_prev[3][139] & 1'b1;
			partial_clause[3][140] 	= partial_clause_prev[3][140] & 1'b1;
			partial_clause[3][141] 	= partial_clause_prev[3][141] & 1'b1;
			partial_clause[3][142] 	= partial_clause_prev[3][142] & 1'b1;
			partial_clause[3][143] 	= partial_clause_prev[3][143] & 1'b1;
			partial_clause[3][144] 	= partial_clause_prev[3][144] & 1'b1;
			partial_clause[3][145] 	= partial_clause_prev[3][145] & 1'b1;
			partial_clause[3][146] 	= partial_clause_prev[3][146] & 1'b1;
			partial_clause[3][147] 	= partial_clause_prev[3][147] & 1'b1;
			partial_clause[3][148] 	= partial_clause_prev[3][148] & 1'b1;
			partial_clause[3][149] 	= partial_clause_prev[3][149] & 1'b1;
			partial_clause[3][150] 	= partial_clause_prev[3][150] & 1'b1;
			partial_clause[3][151] 	= partial_clause_prev[3][151] & 1'b1;
			partial_clause[3][152] 	= partial_clause_prev[3][152] & 1'b1;
			partial_clause[3][153] 	= partial_clause_prev[3][153] & 1'b1;
			partial_clause[3][154] 	= partial_clause_prev[3][154] & 1'b1;
			partial_clause[3][155] 	= partial_clause_prev[3][155] & 1'b1;
			partial_clause[3][156] 	= partial_clause_prev[3][156] & 1'b1;
			partial_clause[3][157] 	= partial_clause_prev[3][157] & 1'b1;
			partial_clause[3][158] 	= partial_clause_prev[3][158] & 1'b1;
			partial_clause[3][159] 	= partial_clause_prev[3][159] & 1'b1;
			partial_clause[3][160] 	= partial_clause_prev[3][160] & 1'b1;
			partial_clause[3][161] 	= partial_clause_prev[3][161] & 1'b1;
			partial_clause[3][162] 	= partial_clause_prev[3][162] & 1'b1;
			partial_clause[3][163] 	= partial_clause_prev[3][163] & 1'b1;
			partial_clause[3][164] 	= partial_clause_prev[3][164] & 1'b1;
			partial_clause[3][165] 	= partial_clause_prev[3][165] & 1'b1;
			partial_clause[3][166] 	= partial_clause_prev[3][166] & 1'b1;
			partial_clause[3][167] 	= partial_clause_prev[3][167] & 1'b1;
			partial_clause[3][168] 	= partial_clause_prev[3][168] & 1'b1;
			partial_clause[3][169] 	= partial_clause_prev[3][169] & 1'b1;
			partial_clause[3][170] 	= partial_clause_prev[3][170] & 1'b1;
			partial_clause[3][171] 	= partial_clause_prev[3][171] & 1'b1;
			partial_clause[3][172] 	= partial_clause_prev[3][172] & 1'b1;
			partial_clause[3][173] 	= partial_clause_prev[3][173] & 1'b1;
			partial_clause[3][174] 	= partial_clause_prev[3][174] & 1'b1;
			partial_clause[3][175] 	= partial_clause_prev[3][175] & 1'b1;
			partial_clause[3][176] 	= partial_clause_prev[3][176] & 1'b1;
			partial_clause[3][177] 	= partial_clause_prev[3][177] & 1'b1;
			partial_clause[3][178] 	= partial_clause_prev[3][178] & 1'b1;
			partial_clause[3][179] 	= partial_clause_prev[3][179] & 1'b1;
			partial_clause[3][180] 	= partial_clause_prev[3][180] & 1'b1;
			partial_clause[3][181] 	= partial_clause_prev[3][181] & 1'b1;
			partial_clause[3][182] 	= partial_clause_prev[3][182] & 1'b1;
			partial_clause[3][183] 	= partial_clause_prev[3][183] & 1'b1;
			partial_clause[3][184] 	= partial_clause_prev[3][184] & 1'b1;
			partial_clause[3][185] 	= partial_clause_prev[3][185] & 1'b1;
			partial_clause[3][186] 	= partial_clause_prev[3][186] & 1'b1;
			partial_clause[3][187] 	= partial_clause_prev[3][187] & 1'b1;
			partial_clause[3][188] 	= partial_clause_prev[3][188] & 1'b1;
			partial_clause[3][189] 	= partial_clause_prev[3][189] & 1'b1;
			partial_clause[3][190] 	= partial_clause_prev[3][190] & 1'b1;
			partial_clause[3][191] 	= partial_clause_prev[3][191] & 1'b1;
			partial_clause[3][192] 	= partial_clause_prev[3][192] & 1'b1;
			partial_clause[3][193] 	= partial_clause_prev[3][193] & 1'b1;
			partial_clause[3][194] 	= partial_clause_prev[3][194] & 1'b1;
			partial_clause[3][195] 	= partial_clause_prev[3][195] & 1'b1;
			partial_clause[3][196] 	= partial_clause_prev[3][196] & 1'b1;
			partial_clause[3][197] 	= partial_clause_prev[3][197] & 1'b1;
			partial_clause[3][198] 	= partial_clause_prev[3][198] & 1'b1;
			partial_clause[3][199] 	= partial_clause_prev[3][199] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & 1'b1;
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & 1'b1;
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & x[12];
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			partial_clause[4][100] 	= partial_clause_prev[4][100] & 1'b1;
			partial_clause[4][101] 	= partial_clause_prev[4][101] & 1'b1;
			partial_clause[4][102] 	= partial_clause_prev[4][102] & 1'b1;
			partial_clause[4][103] 	= partial_clause_prev[4][103] & 1'b1;
			partial_clause[4][104] 	= partial_clause_prev[4][104] & 1'b1;
			partial_clause[4][105] 	= partial_clause_prev[4][105] & 1'b1;
			partial_clause[4][106] 	= partial_clause_prev[4][106] & 1'b1;
			partial_clause[4][107] 	= partial_clause_prev[4][107] & 1'b1;
			partial_clause[4][108] 	= partial_clause_prev[4][108] & 1'b1;
			partial_clause[4][109] 	= partial_clause_prev[4][109] & 1'b1;
			partial_clause[4][110] 	= partial_clause_prev[4][110] & 1'b1;
			partial_clause[4][111] 	= partial_clause_prev[4][111] & 1'b1;
			partial_clause[4][112] 	= partial_clause_prev[4][112] & 1'b1;
			partial_clause[4][113] 	= partial_clause_prev[4][113] & 1'b1;
			partial_clause[4][114] 	= partial_clause_prev[4][114] & 1'b1;
			partial_clause[4][115] 	= partial_clause_prev[4][115] & 1'b1;
			partial_clause[4][116] 	= partial_clause_prev[4][116] & 1'b1;
			partial_clause[4][117] 	= partial_clause_prev[4][117] & 1'b1;
			partial_clause[4][118] 	= partial_clause_prev[4][118] & 1'b1;
			partial_clause[4][119] 	= partial_clause_prev[4][119] & 1'b1;
			partial_clause[4][120] 	= partial_clause_prev[4][120] & 1'b1;
			partial_clause[4][121] 	= partial_clause_prev[4][121] & 1'b1;
			partial_clause[4][122] 	= partial_clause_prev[4][122] & 1'b1;
			partial_clause[4][123] 	= partial_clause_prev[4][123] & 1'b1;
			partial_clause[4][124] 	= partial_clause_prev[4][124] & 1'b1;
			partial_clause[4][125] 	= partial_clause_prev[4][125] & 1'b1;
			partial_clause[4][126] 	= partial_clause_prev[4][126] & 1'b1;
			partial_clause[4][127] 	= partial_clause_prev[4][127] & 1'b1;
			partial_clause[4][128] 	= partial_clause_prev[4][128] & 1'b1;
			partial_clause[4][129] 	= partial_clause_prev[4][129] & 1'b1;
			partial_clause[4][130] 	= partial_clause_prev[4][130] & 1'b1;
			partial_clause[4][131] 	= partial_clause_prev[4][131] & 1'b1;
			partial_clause[4][132] 	= partial_clause_prev[4][132] & 1'b1;
			partial_clause[4][133] 	= partial_clause_prev[4][133] & 1'b1;
			partial_clause[4][134] 	= partial_clause_prev[4][134] & 1'b1;
			partial_clause[4][135] 	= partial_clause_prev[4][135] & 1'b1;
			partial_clause[4][136] 	= partial_clause_prev[4][136] & 1'b1;
			partial_clause[4][137] 	= partial_clause_prev[4][137] & 1'b1;
			partial_clause[4][138] 	= partial_clause_prev[4][138] & 1'b1;
			partial_clause[4][139] 	= partial_clause_prev[4][139] & 1'b1;
			partial_clause[4][140] 	= partial_clause_prev[4][140] & 1'b1;
			partial_clause[4][141] 	= partial_clause_prev[4][141] & 1'b1;
			partial_clause[4][142] 	= partial_clause_prev[4][142] & 1'b1;
			partial_clause[4][143] 	= partial_clause_prev[4][143] & 1'b1;
			partial_clause[4][144] 	= partial_clause_prev[4][144] & 1'b1;
			partial_clause[4][145] 	= partial_clause_prev[4][145] & 1'b1;
			partial_clause[4][146] 	= partial_clause_prev[4][146] & 1'b1;
			partial_clause[4][147] 	= partial_clause_prev[4][147] & 1'b1;
			partial_clause[4][148] 	= partial_clause_prev[4][148] & 1'b1;
			partial_clause[4][149] 	= partial_clause_prev[4][149] & 1'b1;
			partial_clause[4][150] 	= partial_clause_prev[4][150] & 1'b1;
			partial_clause[4][151] 	= partial_clause_prev[4][151] & 1'b1;
			partial_clause[4][152] 	= partial_clause_prev[4][152] & 1'b1;
			partial_clause[4][153] 	= partial_clause_prev[4][153] & 1'b1;
			partial_clause[4][154] 	= partial_clause_prev[4][154] & 1'b1;
			partial_clause[4][155] 	= partial_clause_prev[4][155] & 1'b1;
			partial_clause[4][156] 	= partial_clause_prev[4][156] & 1'b1;
			partial_clause[4][157] 	= partial_clause_prev[4][157] & 1'b1;
			partial_clause[4][158] 	= partial_clause_prev[4][158] & 1'b1;
			partial_clause[4][159] 	= partial_clause_prev[4][159] & 1'b1;
			partial_clause[4][160] 	= partial_clause_prev[4][160] & 1'b1;
			partial_clause[4][161] 	= partial_clause_prev[4][161] & 1'b1;
			partial_clause[4][162] 	= partial_clause_prev[4][162] & 1'b1;
			partial_clause[4][163] 	= partial_clause_prev[4][163] & 1'b1;
			partial_clause[4][164] 	= partial_clause_prev[4][164] & 1'b1;
			partial_clause[4][165] 	= partial_clause_prev[4][165] & 1'b1;
			partial_clause[4][166] 	= partial_clause_prev[4][166] & 1'b1;
			partial_clause[4][167] 	= partial_clause_prev[4][167] & 1'b1;
			partial_clause[4][168] 	= partial_clause_prev[4][168] & 1'b1;
			partial_clause[4][169] 	= partial_clause_prev[4][169] & 1'b1;
			partial_clause[4][170] 	= partial_clause_prev[4][170] & 1'b1;
			partial_clause[4][171] 	= partial_clause_prev[4][171] & 1'b1;
			partial_clause[4][172] 	= partial_clause_prev[4][172] & 1'b1;
			partial_clause[4][173] 	= partial_clause_prev[4][173] & 1'b1;
			partial_clause[4][174] 	= partial_clause_prev[4][174] & 1'b1;
			partial_clause[4][175] 	= partial_clause_prev[4][175] & 1'b1;
			partial_clause[4][176] 	= partial_clause_prev[4][176] & 1'b1;
			partial_clause[4][177] 	= partial_clause_prev[4][177] & 1'b1;
			partial_clause[4][178] 	= partial_clause_prev[4][178] & 1'b1;
			partial_clause[4][179] 	= partial_clause_prev[4][179] & 1'b1;
			partial_clause[4][180] 	= partial_clause_prev[4][180] & 1'b1;
			partial_clause[4][181] 	= partial_clause_prev[4][181] & 1'b1;
			partial_clause[4][182] 	= partial_clause_prev[4][182] & 1'b1;
			partial_clause[4][183] 	= partial_clause_prev[4][183] & 1'b1;
			partial_clause[4][184] 	= partial_clause_prev[4][184] & 1'b1;
			partial_clause[4][185] 	= partial_clause_prev[4][185] & 1'b1;
			partial_clause[4][186] 	= partial_clause_prev[4][186] & 1'b1;
			partial_clause[4][187] 	= partial_clause_prev[4][187] & 1'b1;
			partial_clause[4][188] 	= partial_clause_prev[4][188] & 1'b1;
			partial_clause[4][189] 	= partial_clause_prev[4][189] & 1'b1;
			partial_clause[4][190] 	= partial_clause_prev[4][190] & 1'b1;
			partial_clause[4][191] 	= partial_clause_prev[4][191] & 1'b1;
			partial_clause[4][192] 	= partial_clause_prev[4][192] & 1'b1;
			partial_clause[4][193] 	= partial_clause_prev[4][193] & 1'b1;
			partial_clause[4][194] 	= partial_clause_prev[4][194] & 1'b1;
			partial_clause[4][195] 	= partial_clause_prev[4][195] & 1'b1;
			partial_clause[4][196] 	= partial_clause_prev[4][196] & 1'b1;
			partial_clause[4][197] 	= partial_clause_prev[4][197] & 1'b1;
			partial_clause[4][198] 	= partial_clause_prev[4][198] & 1'b1;
			partial_clause[4][199] 	= partial_clause_prev[4][199] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			partial_clause[5][100] 	= partial_clause_prev[5][100] & 1'b1;
			partial_clause[5][101] 	= partial_clause_prev[5][101] & 1'b1;
			partial_clause[5][102] 	= partial_clause_prev[5][102] & 1'b1;
			partial_clause[5][103] 	= partial_clause_prev[5][103] & 1'b1;
			partial_clause[5][104] 	= partial_clause_prev[5][104] & 1'b1;
			partial_clause[5][105] 	= partial_clause_prev[5][105] & 1'b1;
			partial_clause[5][106] 	= partial_clause_prev[5][106] & 1'b1;
			partial_clause[5][107] 	= partial_clause_prev[5][107] & 1'b1;
			partial_clause[5][108] 	= partial_clause_prev[5][108] & 1'b1;
			partial_clause[5][109] 	= partial_clause_prev[5][109] & 1'b1;
			partial_clause[5][110] 	= partial_clause_prev[5][110] & 1'b1;
			partial_clause[5][111] 	= partial_clause_prev[5][111] & 1'b1;
			partial_clause[5][112] 	= partial_clause_prev[5][112] & 1'b1;
			partial_clause[5][113] 	= partial_clause_prev[5][113] & 1'b1;
			partial_clause[5][114] 	= partial_clause_prev[5][114] & 1'b1;
			partial_clause[5][115] 	= partial_clause_prev[5][115] & 1'b1;
			partial_clause[5][116] 	= partial_clause_prev[5][116] & 1'b1;
			partial_clause[5][117] 	= partial_clause_prev[5][117] & 1'b1;
			partial_clause[5][118] 	= partial_clause_prev[5][118] & 1'b1;
			partial_clause[5][119] 	= partial_clause_prev[5][119] & 1'b1;
			partial_clause[5][120] 	= partial_clause_prev[5][120] & 1'b1;
			partial_clause[5][121] 	= partial_clause_prev[5][121] & 1'b1;
			partial_clause[5][122] 	= partial_clause_prev[5][122] & 1'b1;
			partial_clause[5][123] 	= partial_clause_prev[5][123] & 1'b1;
			partial_clause[5][124] 	= partial_clause_prev[5][124] & 1'b1;
			partial_clause[5][125] 	= partial_clause_prev[5][125] & 1'b1;
			partial_clause[5][126] 	= partial_clause_prev[5][126] & 1'b1;
			partial_clause[5][127] 	= partial_clause_prev[5][127] & 1'b1;
			partial_clause[5][128] 	= partial_clause_prev[5][128] & 1'b1;
			partial_clause[5][129] 	= partial_clause_prev[5][129] & 1'b1;
			partial_clause[5][130] 	= partial_clause_prev[5][130] & 1'b1;
			partial_clause[5][131] 	= partial_clause_prev[5][131] & 1'b1;
			partial_clause[5][132] 	= partial_clause_prev[5][132] & 1'b1;
			partial_clause[5][133] 	= partial_clause_prev[5][133] & 1'b1;
			partial_clause[5][134] 	= partial_clause_prev[5][134] & 1'b1;
			partial_clause[5][135] 	= partial_clause_prev[5][135] & 1'b1;
			partial_clause[5][136] 	= partial_clause_prev[5][136] & 1'b1;
			partial_clause[5][137] 	= partial_clause_prev[5][137] & 1'b1;
			partial_clause[5][138] 	= partial_clause_prev[5][138] & 1'b1;
			partial_clause[5][139] 	= partial_clause_prev[5][139] & 1'b1;
			partial_clause[5][140] 	= partial_clause_prev[5][140] & 1'b1;
			partial_clause[5][141] 	= partial_clause_prev[5][141] & 1'b1;
			partial_clause[5][142] 	= partial_clause_prev[5][142] & 1'b1;
			partial_clause[5][143] 	= partial_clause_prev[5][143] & 1'b1;
			partial_clause[5][144] 	= partial_clause_prev[5][144] & 1'b1;
			partial_clause[5][145] 	= partial_clause_prev[5][145] & 1'b1;
			partial_clause[5][146] 	= partial_clause_prev[5][146] & 1'b1;
			partial_clause[5][147] 	= partial_clause_prev[5][147] & 1'b1;
			partial_clause[5][148] 	= partial_clause_prev[5][148] & 1'b1;
			partial_clause[5][149] 	= partial_clause_prev[5][149] & 1'b1;
			partial_clause[5][150] 	= partial_clause_prev[5][150] & 1'b1;
			partial_clause[5][151] 	= partial_clause_prev[5][151] & 1'b1;
			partial_clause[5][152] 	= partial_clause_prev[5][152] & 1'b1;
			partial_clause[5][153] 	= partial_clause_prev[5][153] & 1'b1;
			partial_clause[5][154] 	= partial_clause_prev[5][154] & 1'b1;
			partial_clause[5][155] 	= partial_clause_prev[5][155] & 1'b1;
			partial_clause[5][156] 	= partial_clause_prev[5][156] & 1'b1;
			partial_clause[5][157] 	= partial_clause_prev[5][157] & 1'b1;
			partial_clause[5][158] 	= partial_clause_prev[5][158] & 1'b1;
			partial_clause[5][159] 	= partial_clause_prev[5][159] & 1'b1;
			partial_clause[5][160] 	= partial_clause_prev[5][160] & 1'b1;
			partial_clause[5][161] 	= partial_clause_prev[5][161] & 1'b1;
			partial_clause[5][162] 	= partial_clause_prev[5][162] & 1'b1;
			partial_clause[5][163] 	= partial_clause_prev[5][163] & 1'b1;
			partial_clause[5][164] 	= partial_clause_prev[5][164] & 1'b1;
			partial_clause[5][165] 	= partial_clause_prev[5][165] & 1'b1;
			partial_clause[5][166] 	= partial_clause_prev[5][166] & 1'b1;
			partial_clause[5][167] 	= partial_clause_prev[5][167] & 1'b1;
			partial_clause[5][168] 	= partial_clause_prev[5][168] & 1'b1;
			partial_clause[5][169] 	= partial_clause_prev[5][169] & 1'b1;
			partial_clause[5][170] 	= partial_clause_prev[5][170] & 1'b1;
			partial_clause[5][171] 	= partial_clause_prev[5][171] & 1'b1;
			partial_clause[5][172] 	= partial_clause_prev[5][172] & 1'b1;
			partial_clause[5][173] 	= partial_clause_prev[5][173] & 1'b1;
			partial_clause[5][174] 	= partial_clause_prev[5][174] & 1'b1;
			partial_clause[5][175] 	= partial_clause_prev[5][175] & 1'b1;
			partial_clause[5][176] 	= partial_clause_prev[5][176] & 1'b1;
			partial_clause[5][177] 	= partial_clause_prev[5][177] & 1'b1;
			partial_clause[5][178] 	= partial_clause_prev[5][178] & 1'b1;
			partial_clause[5][179] 	= partial_clause_prev[5][179] & 1'b1;
			partial_clause[5][180] 	= partial_clause_prev[5][180] & 1'b1;
			partial_clause[5][181] 	= partial_clause_prev[5][181] & 1'b1;
			partial_clause[5][182] 	= partial_clause_prev[5][182] & 1'b1;
			partial_clause[5][183] 	= partial_clause_prev[5][183] & 1'b1;
			partial_clause[5][184] 	= partial_clause_prev[5][184] & 1'b1;
			partial_clause[5][185] 	= partial_clause_prev[5][185] & 1'b1;
			partial_clause[5][186] 	= partial_clause_prev[5][186] & 1'b1;
			partial_clause[5][187] 	= partial_clause_prev[5][187] & 1'b1;
			partial_clause[5][188] 	= partial_clause_prev[5][188] & 1'b1;
			partial_clause[5][189] 	= partial_clause_prev[5][189] & 1'b1;
			partial_clause[5][190] 	= partial_clause_prev[5][190] & 1'b1;
			partial_clause[5][191] 	= partial_clause_prev[5][191] & 1'b1;
			partial_clause[5][192] 	= partial_clause_prev[5][192] & 1'b1;
			partial_clause[5][193] 	= partial_clause_prev[5][193] & 1'b1;
			partial_clause[5][194] 	= partial_clause_prev[5][194] & 1'b1;
			partial_clause[5][195] 	= partial_clause_prev[5][195] & 1'b1;
			partial_clause[5][196] 	= partial_clause_prev[5][196] & 1'b1;
			partial_clause[5][197] 	= partial_clause_prev[5][197] & 1'b1;
			partial_clause[5][198] 	= partial_clause_prev[5][198] & 1'b1;
			partial_clause[5][199] 	= partial_clause_prev[5][199] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & x[6];
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			partial_clause[6][100] 	= partial_clause_prev[6][100] & 1'b1;
			partial_clause[6][101] 	= partial_clause_prev[6][101] & 1'b1;
			partial_clause[6][102] 	= partial_clause_prev[6][102] & 1'b1;
			partial_clause[6][103] 	= partial_clause_prev[6][103] & 1'b1;
			partial_clause[6][104] 	= partial_clause_prev[6][104] & 1'b1;
			partial_clause[6][105] 	= partial_clause_prev[6][105] & 1'b1;
			partial_clause[6][106] 	= partial_clause_prev[6][106] & 1'b1;
			partial_clause[6][107] 	= partial_clause_prev[6][107] & 1'b1;
			partial_clause[6][108] 	= partial_clause_prev[6][108] & 1'b1;
			partial_clause[6][109] 	= partial_clause_prev[6][109] & 1'b1;
			partial_clause[6][110] 	= partial_clause_prev[6][110] & 1'b1;
			partial_clause[6][111] 	= partial_clause_prev[6][111] & 1'b1;
			partial_clause[6][112] 	= partial_clause_prev[6][112] & 1'b1;
			partial_clause[6][113] 	= partial_clause_prev[6][113] & 1'b1;
			partial_clause[6][114] 	= partial_clause_prev[6][114] & 1'b1;
			partial_clause[6][115] 	= partial_clause_prev[6][115] & 1'b1;
			partial_clause[6][116] 	= partial_clause_prev[6][116] & 1'b1;
			partial_clause[6][117] 	= partial_clause_prev[6][117] & 1'b1;
			partial_clause[6][118] 	= partial_clause_prev[6][118] & 1'b1;
			partial_clause[6][119] 	= partial_clause_prev[6][119] & 1'b1;
			partial_clause[6][120] 	= partial_clause_prev[6][120] & 1'b1;
			partial_clause[6][121] 	= partial_clause_prev[6][121] & 1'b1;
			partial_clause[6][122] 	= partial_clause_prev[6][122] & 1'b1;
			partial_clause[6][123] 	= partial_clause_prev[6][123] & 1'b1;
			partial_clause[6][124] 	= partial_clause_prev[6][124] & 1'b1;
			partial_clause[6][125] 	= partial_clause_prev[6][125] & 1'b1;
			partial_clause[6][126] 	= partial_clause_prev[6][126] & 1'b1;
			partial_clause[6][127] 	= partial_clause_prev[6][127] & 1'b1;
			partial_clause[6][128] 	= partial_clause_prev[6][128] & 1'b1;
			partial_clause[6][129] 	= partial_clause_prev[6][129] & 1'b1;
			partial_clause[6][130] 	= partial_clause_prev[6][130] & 1'b1;
			partial_clause[6][131] 	= partial_clause_prev[6][131] & 1'b1;
			partial_clause[6][132] 	= partial_clause_prev[6][132] & 1'b1;
			partial_clause[6][133] 	= partial_clause_prev[6][133] & 1'b1;
			partial_clause[6][134] 	= partial_clause_prev[6][134] & 1'b1;
			partial_clause[6][135] 	= partial_clause_prev[6][135] & 1'b1;
			partial_clause[6][136] 	= partial_clause_prev[6][136] & 1'b1;
			partial_clause[6][137] 	= partial_clause_prev[6][137] & 1'b1;
			partial_clause[6][138] 	= partial_clause_prev[6][138] & 1'b1;
			partial_clause[6][139] 	= partial_clause_prev[6][139] & 1'b1;
			partial_clause[6][140] 	= partial_clause_prev[6][140] & 1'b1;
			partial_clause[6][141] 	= partial_clause_prev[6][141] & 1'b1;
			partial_clause[6][142] 	= partial_clause_prev[6][142] & 1'b1;
			partial_clause[6][143] 	= partial_clause_prev[6][143] & 1'b1;
			partial_clause[6][144] 	= partial_clause_prev[6][144] & 1'b1;
			partial_clause[6][145] 	= partial_clause_prev[6][145] & 1'b1;
			partial_clause[6][146] 	= partial_clause_prev[6][146] & 1'b1;
			partial_clause[6][147] 	= partial_clause_prev[6][147] & 1'b1;
			partial_clause[6][148] 	= partial_clause_prev[6][148] & 1'b1;
			partial_clause[6][149] 	= partial_clause_prev[6][149] & 1'b1;
			partial_clause[6][150] 	= partial_clause_prev[6][150] & 1'b1;
			partial_clause[6][151] 	= partial_clause_prev[6][151] & 1'b1;
			partial_clause[6][152] 	= partial_clause_prev[6][152] & 1'b1;
			partial_clause[6][153] 	= partial_clause_prev[6][153] & 1'b1;
			partial_clause[6][154] 	= partial_clause_prev[6][154] & 1'b1;
			partial_clause[6][155] 	= partial_clause_prev[6][155] & 1'b1;
			partial_clause[6][156] 	= partial_clause_prev[6][156] & 1'b1;
			partial_clause[6][157] 	= partial_clause_prev[6][157] & 1'b1;
			partial_clause[6][158] 	= partial_clause_prev[6][158] & 1'b1;
			partial_clause[6][159] 	= partial_clause_prev[6][159] & 1'b1;
			partial_clause[6][160] 	= partial_clause_prev[6][160] & 1'b1;
			partial_clause[6][161] 	= partial_clause_prev[6][161] & 1'b1;
			partial_clause[6][162] 	= partial_clause_prev[6][162] & 1'b1;
			partial_clause[6][163] 	= partial_clause_prev[6][163] & 1'b1;
			partial_clause[6][164] 	= partial_clause_prev[6][164] & 1'b1;
			partial_clause[6][165] 	= partial_clause_prev[6][165] & 1'b1;
			partial_clause[6][166] 	= partial_clause_prev[6][166] & 1'b1;
			partial_clause[6][167] 	= partial_clause_prev[6][167] & 1'b1;
			partial_clause[6][168] 	= partial_clause_prev[6][168] & 1'b1;
			partial_clause[6][169] 	= partial_clause_prev[6][169] & 1'b1;
			partial_clause[6][170] 	= partial_clause_prev[6][170] & 1'b1;
			partial_clause[6][171] 	= partial_clause_prev[6][171] & 1'b1;
			partial_clause[6][172] 	= partial_clause_prev[6][172] & 1'b1;
			partial_clause[6][173] 	= partial_clause_prev[6][173] & 1'b1;
			partial_clause[6][174] 	= partial_clause_prev[6][174] & 1'b1;
			partial_clause[6][175] 	= partial_clause_prev[6][175] & 1'b1;
			partial_clause[6][176] 	= partial_clause_prev[6][176] & 1'b1;
			partial_clause[6][177] 	= partial_clause_prev[6][177] & 1'b1;
			partial_clause[6][178] 	= partial_clause_prev[6][178] & 1'b1;
			partial_clause[6][179] 	= partial_clause_prev[6][179] & 1'b1;
			partial_clause[6][180] 	= partial_clause_prev[6][180] & 1'b1;
			partial_clause[6][181] 	= partial_clause_prev[6][181] & 1'b1;
			partial_clause[6][182] 	= partial_clause_prev[6][182] & 1'b1;
			partial_clause[6][183] 	= partial_clause_prev[6][183] & 1'b1;
			partial_clause[6][184] 	= partial_clause_prev[6][184] & 1'b1;
			partial_clause[6][185] 	= partial_clause_prev[6][185] & 1'b1;
			partial_clause[6][186] 	= partial_clause_prev[6][186] & 1'b1;
			partial_clause[6][187] 	= partial_clause_prev[6][187] & ~x[7];
			partial_clause[6][188] 	= partial_clause_prev[6][188] & 1'b1;
			partial_clause[6][189] 	= partial_clause_prev[6][189] & 1'b1;
			partial_clause[6][190] 	= partial_clause_prev[6][190] & 1'b1;
			partial_clause[6][191] 	= partial_clause_prev[6][191] & 1'b1;
			partial_clause[6][192] 	= partial_clause_prev[6][192] & 1'b1;
			partial_clause[6][193] 	= partial_clause_prev[6][193] & 1'b1;
			partial_clause[6][194] 	= partial_clause_prev[6][194] & 1'b1;
			partial_clause[6][195] 	= partial_clause_prev[6][195] & 1'b1;
			partial_clause[6][196] 	= partial_clause_prev[6][196] & 1'b1;
			partial_clause[6][197] 	= partial_clause_prev[6][197] & 1'b1;
			partial_clause[6][198] 	= partial_clause_prev[6][198] & 1'b1;
			partial_clause[6][199] 	= partial_clause_prev[6][199] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & x[5];
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			partial_clause[7][100] 	= partial_clause_prev[7][100] & 1'b1;
			partial_clause[7][101] 	= partial_clause_prev[7][101] & 1'b1;
			partial_clause[7][102] 	= partial_clause_prev[7][102] & 1'b1;
			partial_clause[7][103] 	= partial_clause_prev[7][103] & 1'b1;
			partial_clause[7][104] 	= partial_clause_prev[7][104] & 1'b1;
			partial_clause[7][105] 	= partial_clause_prev[7][105] & 1'b1;
			partial_clause[7][106] 	= partial_clause_prev[7][106] & 1'b1;
			partial_clause[7][107] 	= partial_clause_prev[7][107] & 1'b1;
			partial_clause[7][108] 	= partial_clause_prev[7][108] & 1'b1;
			partial_clause[7][109] 	= partial_clause_prev[7][109] & 1'b1;
			partial_clause[7][110] 	= partial_clause_prev[7][110] & 1'b1;
			partial_clause[7][111] 	= partial_clause_prev[7][111] & 1'b1;
			partial_clause[7][112] 	= partial_clause_prev[7][112] & 1'b1;
			partial_clause[7][113] 	= partial_clause_prev[7][113] & 1'b1;
			partial_clause[7][114] 	= partial_clause_prev[7][114] & 1'b1;
			partial_clause[7][115] 	= partial_clause_prev[7][115] & 1'b1;
			partial_clause[7][116] 	= partial_clause_prev[7][116] & 1'b1;
			partial_clause[7][117] 	= partial_clause_prev[7][117] & 1'b1;
			partial_clause[7][118] 	= partial_clause_prev[7][118] & 1'b1;
			partial_clause[7][119] 	= partial_clause_prev[7][119] & 1'b1;
			partial_clause[7][120] 	= partial_clause_prev[7][120] & 1'b1;
			partial_clause[7][121] 	= partial_clause_prev[7][121] & 1'b1;
			partial_clause[7][122] 	= partial_clause_prev[7][122] & 1'b1;
			partial_clause[7][123] 	= partial_clause_prev[7][123] & 1'b1;
			partial_clause[7][124] 	= partial_clause_prev[7][124] & 1'b1;
			partial_clause[7][125] 	= partial_clause_prev[7][125] & 1'b1;
			partial_clause[7][126] 	= partial_clause_prev[7][126] & 1'b1;
			partial_clause[7][127] 	= partial_clause_prev[7][127] & 1'b1;
			partial_clause[7][128] 	= partial_clause_prev[7][128] & 1'b1;
			partial_clause[7][129] 	= partial_clause_prev[7][129] & 1'b1;
			partial_clause[7][130] 	= partial_clause_prev[7][130] & ~x[1];
			partial_clause[7][131] 	= partial_clause_prev[7][131] & 1'b1;
			partial_clause[7][132] 	= partial_clause_prev[7][132] & 1'b1;
			partial_clause[7][133] 	= partial_clause_prev[7][133] & 1'b1;
			partial_clause[7][134] 	= partial_clause_prev[7][134] & 1'b1;
			partial_clause[7][135] 	= partial_clause_prev[7][135] & 1'b1;
			partial_clause[7][136] 	= partial_clause_prev[7][136] & 1'b1;
			partial_clause[7][137] 	= partial_clause_prev[7][137] & 1'b1;
			partial_clause[7][138] 	= partial_clause_prev[7][138] & 1'b1;
			partial_clause[7][139] 	= partial_clause_prev[7][139] & 1'b1;
			partial_clause[7][140] 	= partial_clause_prev[7][140] & 1'b1;
			partial_clause[7][141] 	= partial_clause_prev[7][141] & 1'b1;
			partial_clause[7][142] 	= partial_clause_prev[7][142] & 1'b1;
			partial_clause[7][143] 	= partial_clause_prev[7][143] & 1'b1;
			partial_clause[7][144] 	= partial_clause_prev[7][144] & 1'b1;
			partial_clause[7][145] 	= partial_clause_prev[7][145] & 1'b1;
			partial_clause[7][146] 	= partial_clause_prev[7][146] & 1'b1;
			partial_clause[7][147] 	= partial_clause_prev[7][147] & 1'b1;
			partial_clause[7][148] 	= partial_clause_prev[7][148] & 1'b1;
			partial_clause[7][149] 	= partial_clause_prev[7][149] & 1'b1;
			partial_clause[7][150] 	= partial_clause_prev[7][150] & 1'b1;
			partial_clause[7][151] 	= partial_clause_prev[7][151] & 1'b1;
			partial_clause[7][152] 	= partial_clause_prev[7][152] & 1'b1;
			partial_clause[7][153] 	= partial_clause_prev[7][153] & 1'b1;
			partial_clause[7][154] 	= partial_clause_prev[7][154] & 1'b1;
			partial_clause[7][155] 	= partial_clause_prev[7][155] & 1'b1;
			partial_clause[7][156] 	= partial_clause_prev[7][156] & 1'b1;
			partial_clause[7][157] 	= partial_clause_prev[7][157] & 1'b1;
			partial_clause[7][158] 	= partial_clause_prev[7][158] & 1'b1;
			partial_clause[7][159] 	= partial_clause_prev[7][159] & 1'b1;
			partial_clause[7][160] 	= partial_clause_prev[7][160] & 1'b1;
			partial_clause[7][161] 	= partial_clause_prev[7][161] & 1'b1;
			partial_clause[7][162] 	= partial_clause_prev[7][162] & 1'b1;
			partial_clause[7][163] 	= partial_clause_prev[7][163] & 1'b1;
			partial_clause[7][164] 	= partial_clause_prev[7][164] & 1'b1;
			partial_clause[7][165] 	= partial_clause_prev[7][165] & 1'b1;
			partial_clause[7][166] 	= partial_clause_prev[7][166] & 1'b1;
			partial_clause[7][167] 	= partial_clause_prev[7][167] & 1'b1;
			partial_clause[7][168] 	= partial_clause_prev[7][168] & 1'b1;
			partial_clause[7][169] 	= partial_clause_prev[7][169] & 1'b1;
			partial_clause[7][170] 	= partial_clause_prev[7][170] & 1'b1;
			partial_clause[7][171] 	= partial_clause_prev[7][171] & 1'b1;
			partial_clause[7][172] 	= partial_clause_prev[7][172] & 1'b1;
			partial_clause[7][173] 	= partial_clause_prev[7][173] & 1'b1;
			partial_clause[7][174] 	= partial_clause_prev[7][174] & 1'b1;
			partial_clause[7][175] 	= partial_clause_prev[7][175] & 1'b1;
			partial_clause[7][176] 	= partial_clause_prev[7][176] & 1'b1;
			partial_clause[7][177] 	= partial_clause_prev[7][177] & 1'b1;
			partial_clause[7][178] 	= partial_clause_prev[7][178] & 1'b1;
			partial_clause[7][179] 	= partial_clause_prev[7][179] & 1'b1;
			partial_clause[7][180] 	= partial_clause_prev[7][180] & 1'b1;
			partial_clause[7][181] 	= partial_clause_prev[7][181] & 1'b1;
			partial_clause[7][182] 	= partial_clause_prev[7][182] & 1'b1;
			partial_clause[7][183] 	= partial_clause_prev[7][183] & 1'b1;
			partial_clause[7][184] 	= partial_clause_prev[7][184] & 1'b1;
			partial_clause[7][185] 	= partial_clause_prev[7][185] & 1'b1;
			partial_clause[7][186] 	= partial_clause_prev[7][186] & 1'b1;
			partial_clause[7][187] 	= partial_clause_prev[7][187] & 1'b1;
			partial_clause[7][188] 	= partial_clause_prev[7][188] & 1'b1;
			partial_clause[7][189] 	= partial_clause_prev[7][189] & 1'b1;
			partial_clause[7][190] 	= partial_clause_prev[7][190] & 1'b1;
			partial_clause[7][191] 	= partial_clause_prev[7][191] & 1'b1;
			partial_clause[7][192] 	= partial_clause_prev[7][192] & 1'b1;
			partial_clause[7][193] 	= partial_clause_prev[7][193] & 1'b1;
			partial_clause[7][194] 	= partial_clause_prev[7][194] & 1'b1;
			partial_clause[7][195] 	= partial_clause_prev[7][195] & 1'b1;
			partial_clause[7][196] 	= partial_clause_prev[7][196] & 1'b1;
			partial_clause[7][197] 	= partial_clause_prev[7][197] & 1'b1;
			partial_clause[7][198] 	= partial_clause_prev[7][198] & 1'b1;
			partial_clause[7][199] 	= partial_clause_prev[7][199] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & ~x[4];
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & x[9];
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & x[6];
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & x[12];
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			partial_clause[8][100] 	= partial_clause_prev[8][100] & 1'b1;
			partial_clause[8][101] 	= partial_clause_prev[8][101] & 1'b1;
			partial_clause[8][102] 	= partial_clause_prev[8][102] & 1'b1;
			partial_clause[8][103] 	= partial_clause_prev[8][103] & 1'b1;
			partial_clause[8][104] 	= partial_clause_prev[8][104] & 1'b1;
			partial_clause[8][105] 	= partial_clause_prev[8][105] & 1'b1;
			partial_clause[8][106] 	= partial_clause_prev[8][106] & 1'b1;
			partial_clause[8][107] 	= partial_clause_prev[8][107] & 1'b1;
			partial_clause[8][108] 	= partial_clause_prev[8][108] & 1'b1;
			partial_clause[8][109] 	= partial_clause_prev[8][109] & 1'b1;
			partial_clause[8][110] 	= partial_clause_prev[8][110] & 1'b1;
			partial_clause[8][111] 	= partial_clause_prev[8][111] & x[0];
			partial_clause[8][112] 	= partial_clause_prev[8][112] & 1'b1;
			partial_clause[8][113] 	= partial_clause_prev[8][113] & 1'b1;
			partial_clause[8][114] 	= partial_clause_prev[8][114] & 1'b1;
			partial_clause[8][115] 	= partial_clause_prev[8][115] & 1'b1;
			partial_clause[8][116] 	= partial_clause_prev[8][116] & 1'b1;
			partial_clause[8][117] 	= partial_clause_prev[8][117] & 1'b1;
			partial_clause[8][118] 	= partial_clause_prev[8][118] & 1'b1;
			partial_clause[8][119] 	= partial_clause_prev[8][119] & 1'b1;
			partial_clause[8][120] 	= partial_clause_prev[8][120] & 1'b1;
			partial_clause[8][121] 	= partial_clause_prev[8][121] & 1'b1;
			partial_clause[8][122] 	= partial_clause_prev[8][122] & 1'b1;
			partial_clause[8][123] 	= partial_clause_prev[8][123] & 1'b1;
			partial_clause[8][124] 	= partial_clause_prev[8][124] & 1'b1;
			partial_clause[8][125] 	= partial_clause_prev[8][125] & 1'b1;
			partial_clause[8][126] 	= partial_clause_prev[8][126] & 1'b1;
			partial_clause[8][127] 	= partial_clause_prev[8][127] & 1'b1;
			partial_clause[8][128] 	= partial_clause_prev[8][128] & 1'b1;
			partial_clause[8][129] 	= partial_clause_prev[8][129] & 1'b1;
			partial_clause[8][130] 	= partial_clause_prev[8][130] & 1'b1;
			partial_clause[8][131] 	= partial_clause_prev[8][131] & 1'b1;
			partial_clause[8][132] 	= partial_clause_prev[8][132] & 1'b1;
			partial_clause[8][133] 	= partial_clause_prev[8][133] & 1'b1;
			partial_clause[8][134] 	= partial_clause_prev[8][134] & 1'b1;
			partial_clause[8][135] 	= partial_clause_prev[8][135] & 1'b1;
			partial_clause[8][136] 	= partial_clause_prev[8][136] & 1'b1;
			partial_clause[8][137] 	= partial_clause_prev[8][137] & 1'b1;
			partial_clause[8][138] 	= partial_clause_prev[8][138] & 1'b1;
			partial_clause[8][139] 	= partial_clause_prev[8][139] & 1'b1;
			partial_clause[8][140] 	= partial_clause_prev[8][140] & 1'b1;
			partial_clause[8][141] 	= partial_clause_prev[8][141] & 1'b1;
			partial_clause[8][142] 	= partial_clause_prev[8][142] & 1'b1;
			partial_clause[8][143] 	= partial_clause_prev[8][143] & 1'b1;
			partial_clause[8][144] 	= partial_clause_prev[8][144] & 1'b1;
			partial_clause[8][145] 	= partial_clause_prev[8][145] & 1'b1;
			partial_clause[8][146] 	= partial_clause_prev[8][146] & 1'b1;
			partial_clause[8][147] 	= partial_clause_prev[8][147] & 1'b1;
			partial_clause[8][148] 	= partial_clause_prev[8][148] & 1'b1;
			partial_clause[8][149] 	= partial_clause_prev[8][149] & 1'b1;
			partial_clause[8][150] 	= partial_clause_prev[8][150] & 1'b1;
			partial_clause[8][151] 	= partial_clause_prev[8][151] & 1'b1;
			partial_clause[8][152] 	= partial_clause_prev[8][152] & 1'b1;
			partial_clause[8][153] 	= partial_clause_prev[8][153] & 1'b1;
			partial_clause[8][154] 	= partial_clause_prev[8][154] & 1'b1;
			partial_clause[8][155] 	= partial_clause_prev[8][155] & 1'b1;
			partial_clause[8][156] 	= partial_clause_prev[8][156] & 1'b1;
			partial_clause[8][157] 	= partial_clause_prev[8][157] & 1'b1;
			partial_clause[8][158] 	= partial_clause_prev[8][158] & 1'b1;
			partial_clause[8][159] 	= partial_clause_prev[8][159] & 1'b1;
			partial_clause[8][160] 	= partial_clause_prev[8][160] & 1'b1;
			partial_clause[8][161] 	= partial_clause_prev[8][161] & 1'b1;
			partial_clause[8][162] 	= partial_clause_prev[8][162] & 1'b1;
			partial_clause[8][163] 	= partial_clause_prev[8][163] & 1'b1;
			partial_clause[8][164] 	= partial_clause_prev[8][164] & 1'b1;
			partial_clause[8][165] 	= partial_clause_prev[8][165] & 1'b1;
			partial_clause[8][166] 	= partial_clause_prev[8][166] & 1'b1;
			partial_clause[8][167] 	= partial_clause_prev[8][167] & 1'b1;
			partial_clause[8][168] 	= partial_clause_prev[8][168] & 1'b1;
			partial_clause[8][169] 	= partial_clause_prev[8][169] & 1'b1;
			partial_clause[8][170] 	= partial_clause_prev[8][170] & 1'b1;
			partial_clause[8][171] 	= partial_clause_prev[8][171] & 1'b1;
			partial_clause[8][172] 	= partial_clause_prev[8][172] & 1'b1;
			partial_clause[8][173] 	= partial_clause_prev[8][173] & 1'b1;
			partial_clause[8][174] 	= partial_clause_prev[8][174] & 1'b1;
			partial_clause[8][175] 	= partial_clause_prev[8][175] & 1'b1;
			partial_clause[8][176] 	= partial_clause_prev[8][176] & 1'b1;
			partial_clause[8][177] 	= partial_clause_prev[8][177] & 1'b1;
			partial_clause[8][178] 	= partial_clause_prev[8][178] & 1'b1;
			partial_clause[8][179] 	= partial_clause_prev[8][179] & 1'b1;
			partial_clause[8][180] 	= partial_clause_prev[8][180] & 1'b1;
			partial_clause[8][181] 	= partial_clause_prev[8][181] & 1'b1;
			partial_clause[8][182] 	= partial_clause_prev[8][182] & 1'b1;
			partial_clause[8][183] 	= partial_clause_prev[8][183] & 1'b1;
			partial_clause[8][184] 	= partial_clause_prev[8][184] & 1'b1;
			partial_clause[8][185] 	= partial_clause_prev[8][185] & 1'b1;
			partial_clause[8][186] 	= partial_clause_prev[8][186] & 1'b1;
			partial_clause[8][187] 	= partial_clause_prev[8][187] & 1'b1;
			partial_clause[8][188] 	= partial_clause_prev[8][188] & 1'b1;
			partial_clause[8][189] 	= partial_clause_prev[8][189] & 1'b1;
			partial_clause[8][190] 	= partial_clause_prev[8][190] & 1'b1;
			partial_clause[8][191] 	= partial_clause_prev[8][191] & 1'b1;
			partial_clause[8][192] 	= partial_clause_prev[8][192] & 1'b1;
			partial_clause[8][193] 	= partial_clause_prev[8][193] & 1'b1;
			partial_clause[8][194] 	= partial_clause_prev[8][194] & 1'b1;
			partial_clause[8][195] 	= partial_clause_prev[8][195] & 1'b1;
			partial_clause[8][196] 	= partial_clause_prev[8][196] & 1'b1;
			partial_clause[8][197] 	= partial_clause_prev[8][197] & 1'b1;
			partial_clause[8][198] 	= partial_clause_prev[8][198] & 1'b1;
			partial_clause[8][199] 	= partial_clause_prev[8][199] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & 1'b1;
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
			partial_clause[9][100] 	= partial_clause_prev[9][100] & 1'b1;
			partial_clause[9][101] 	= partial_clause_prev[9][101] & 1'b1;
			partial_clause[9][102] 	= partial_clause_prev[9][102] & 1'b1;
			partial_clause[9][103] 	= partial_clause_prev[9][103] & 1'b1;
			partial_clause[9][104] 	= partial_clause_prev[9][104] & 1'b1;
			partial_clause[9][105] 	= partial_clause_prev[9][105] & 1'b1;
			partial_clause[9][106] 	= partial_clause_prev[9][106] & 1'b1;
			partial_clause[9][107] 	= partial_clause_prev[9][107] & 1'b1;
			partial_clause[9][108] 	= partial_clause_prev[9][108] & 1'b1;
			partial_clause[9][109] 	= partial_clause_prev[9][109] & 1'b1;
			partial_clause[9][110] 	= partial_clause_prev[9][110] & 1'b1;
			partial_clause[9][111] 	= partial_clause_prev[9][111] & 1'b1;
			partial_clause[9][112] 	= partial_clause_prev[9][112] & 1'b1;
			partial_clause[9][113] 	= partial_clause_prev[9][113] & 1'b1;
			partial_clause[9][114] 	= partial_clause_prev[9][114] & 1'b1;
			partial_clause[9][115] 	= partial_clause_prev[9][115] & 1'b1;
			partial_clause[9][116] 	= partial_clause_prev[9][116] & 1'b1;
			partial_clause[9][117] 	= partial_clause_prev[9][117] & 1'b1;
			partial_clause[9][118] 	= partial_clause_prev[9][118] & 1'b1;
			partial_clause[9][119] 	= partial_clause_prev[9][119] & 1'b1;
			partial_clause[9][120] 	= partial_clause_prev[9][120] & 1'b1;
			partial_clause[9][121] 	= partial_clause_prev[9][121] & 1'b1;
			partial_clause[9][122] 	= partial_clause_prev[9][122] & 1'b1;
			partial_clause[9][123] 	= partial_clause_prev[9][123] & 1'b1;
			partial_clause[9][124] 	= partial_clause_prev[9][124] & 1'b1;
			partial_clause[9][125] 	= partial_clause_prev[9][125] & 1'b1;
			partial_clause[9][126] 	= partial_clause_prev[9][126] & 1'b1;
			partial_clause[9][127] 	= partial_clause_prev[9][127] & 1'b1;
			partial_clause[9][128] 	= partial_clause_prev[9][128] & 1'b1;
			partial_clause[9][129] 	= partial_clause_prev[9][129] & 1'b1;
			partial_clause[9][130] 	= partial_clause_prev[9][130] & 1'b1;
			partial_clause[9][131] 	= partial_clause_prev[9][131] & 1'b1;
			partial_clause[9][132] 	= partial_clause_prev[9][132] & 1'b1;
			partial_clause[9][133] 	= partial_clause_prev[9][133] & 1'b1;
			partial_clause[9][134] 	= partial_clause_prev[9][134] & 1'b1;
			partial_clause[9][135] 	= partial_clause_prev[9][135] & 1'b1;
			partial_clause[9][136] 	= partial_clause_prev[9][136] & 1'b1;
			partial_clause[9][137] 	= partial_clause_prev[9][137] & 1'b1;
			partial_clause[9][138] 	= partial_clause_prev[9][138] & 1'b1;
			partial_clause[9][139] 	= partial_clause_prev[9][139] & 1'b1;
			partial_clause[9][140] 	= partial_clause_prev[9][140] & 1'b1;
			partial_clause[9][141] 	= partial_clause_prev[9][141] & 1'b1;
			partial_clause[9][142] 	= partial_clause_prev[9][142] & 1'b1;
			partial_clause[9][143] 	= partial_clause_prev[9][143] & 1'b1;
			partial_clause[9][144] 	= partial_clause_prev[9][144] & 1'b1;
			partial_clause[9][145] 	= partial_clause_prev[9][145] & 1'b1;
			partial_clause[9][146] 	= partial_clause_prev[9][146] & 1'b1;
			partial_clause[9][147] 	= partial_clause_prev[9][147] & 1'b1;
			partial_clause[9][148] 	= partial_clause_prev[9][148] & 1'b1;
			partial_clause[9][149] 	= partial_clause_prev[9][149] & 1'b1;
			partial_clause[9][150] 	= partial_clause_prev[9][150] & 1'b1;
			partial_clause[9][151] 	= partial_clause_prev[9][151] & 1'b1;
			partial_clause[9][152] 	= partial_clause_prev[9][152] & 1'b1;
			partial_clause[9][153] 	= partial_clause_prev[9][153] & 1'b1;
			partial_clause[9][154] 	= partial_clause_prev[9][154] & 1'b1;
			partial_clause[9][155] 	= partial_clause_prev[9][155] & 1'b1;
			partial_clause[9][156] 	= partial_clause_prev[9][156] & 1'b1;
			partial_clause[9][157] 	= partial_clause_prev[9][157] & 1'b1;
			partial_clause[9][158] 	= partial_clause_prev[9][158] & 1'b1;
			partial_clause[9][159] 	= partial_clause_prev[9][159] & 1'b1;
			partial_clause[9][160] 	= partial_clause_prev[9][160] & 1'b1;
			partial_clause[9][161] 	= partial_clause_prev[9][161] & 1'b1;
			partial_clause[9][162] 	= partial_clause_prev[9][162] & 1'b1;
			partial_clause[9][163] 	= partial_clause_prev[9][163] & 1'b1;
			partial_clause[9][164] 	= partial_clause_prev[9][164] & 1'b1;
			partial_clause[9][165] 	= partial_clause_prev[9][165] & 1'b1;
			partial_clause[9][166] 	= partial_clause_prev[9][166] & 1'b1;
			partial_clause[9][167] 	= partial_clause_prev[9][167] & 1'b1;
			partial_clause[9][168] 	= partial_clause_prev[9][168] & 1'b1;
			partial_clause[9][169] 	= partial_clause_prev[9][169] & 1'b1;
			partial_clause[9][170] 	= partial_clause_prev[9][170] & 1'b1;
			partial_clause[9][171] 	= partial_clause_prev[9][171] & 1'b1;
			partial_clause[9][172] 	= partial_clause_prev[9][172] & 1'b1;
			partial_clause[9][173] 	= partial_clause_prev[9][173] & 1'b1;
			partial_clause[9][174] 	= partial_clause_prev[9][174] & 1'b1;
			partial_clause[9][175] 	= partial_clause_prev[9][175] & 1'b1;
			partial_clause[9][176] 	= partial_clause_prev[9][176] & 1'b1;
			partial_clause[9][177] 	= partial_clause_prev[9][177] & 1'b1;
			partial_clause[9][178] 	= partial_clause_prev[9][178] & 1'b1;
			partial_clause[9][179] 	= partial_clause_prev[9][179] & 1'b1;
			partial_clause[9][180] 	= partial_clause_prev[9][180] & 1'b1;
			partial_clause[9][181] 	= partial_clause_prev[9][181] & 1'b1;
			partial_clause[9][182] 	= partial_clause_prev[9][182] & 1'b1;
			partial_clause[9][183] 	= partial_clause_prev[9][183] & 1'b1;
			partial_clause[9][184] 	= partial_clause_prev[9][184] & 1'b1;
			partial_clause[9][185] 	= partial_clause_prev[9][185] & 1'b1;
			partial_clause[9][186] 	= partial_clause_prev[9][186] & 1'b1;
			partial_clause[9][187] 	= partial_clause_prev[9][187] & 1'b1;
			partial_clause[9][188] 	= partial_clause_prev[9][188] & 1'b1;
			partial_clause[9][189] 	= partial_clause_prev[9][189] & 1'b1;
			partial_clause[9][190] 	= partial_clause_prev[9][190] & 1'b1;
			partial_clause[9][191] 	= partial_clause_prev[9][191] & 1'b1;
			partial_clause[9][192] 	= partial_clause_prev[9][192] & 1'b1;
			partial_clause[9][193] 	= partial_clause_prev[9][193] & 1'b1;
			partial_clause[9][194] 	= partial_clause_prev[9][194] & 1'b1;
			partial_clause[9][195] 	= partial_clause_prev[9][195] & 1'b1;
			partial_clause[9][196] 	= partial_clause_prev[9][196] & 1'b1;
			partial_clause[9][197] 	= partial_clause_prev[9][197] & 1'b1;
			partial_clause[9][198] 	= partial_clause_prev[9][198] & 1'b1;
			partial_clause[9][199] 	= partial_clause_prev[9][199] & 1'b1;
		end
	end
endmodule


