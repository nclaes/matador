module HCB_0 (x, partial_clause, clk, valid);
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= 1'b1;
			partial_clause[0][1] 	= ~x[31];
			partial_clause[0][2] 	= 1'b1;
			partial_clause[0][3] 	= ~x[33];
			partial_clause[0][4] 	= 1'b1;
			partial_clause[0][5] 	= 1'b1;
			partial_clause[0][6] 	= ~x[29];
			partial_clause[0][7] 	= ~x[0] & ~x[53];
			partial_clause[0][8] 	= ~x[11];
			partial_clause[0][9] 	= 1'b1;
			partial_clause[0][10] 	= 1'b1;
			partial_clause[0][11] 	= 1'b1;
			partial_clause[0][12] 	= 1'b1;
			partial_clause[0][13] 	= 1'b1;
			partial_clause[0][14] 	= 1'b1;
			partial_clause[0][15] 	= ~x[32];
			partial_clause[0][16] 	= 1'b1;
			partial_clause[0][17] 	= ~x[30] & ~x[59];
			partial_clause[0][18] 	= 1'b1;
			partial_clause[0][19] 	= 1'b1;
			partial_clause[0][20] 	= 1'b1;
			partial_clause[0][21] 	= 1'b1;
			partial_clause[0][22] 	= 1'b1;
			partial_clause[0][23] 	= ~x[30];
			partial_clause[0][24] 	= ~x[56];
			partial_clause[0][25] 	= 1'b1;
			partial_clause[0][26] 	= 1'b1;
			partial_clause[0][27] 	= ~x[33];
			partial_clause[0][28] 	= ~x[58];
			partial_clause[0][29] 	= 1'b1;
			partial_clause[0][30] 	= ~x[55];
			partial_clause[0][31] 	= 1'b1;
			partial_clause[0][32] 	= 1'b1;
			partial_clause[0][33] 	= 1'b1;
			partial_clause[0][34] 	= ~x[16];
			partial_clause[0][35] 	= 1'b1;
			partial_clause[0][36] 	= 1'b1;
			partial_clause[0][37] 	= 1'b1;
			partial_clause[0][38] 	= 1'b1;
			partial_clause[0][39] 	= 1'b1;
			partial_clause[0][40] 	= 1'b1;
			partial_clause[0][41] 	= ~x[47];
			partial_clause[0][42] 	= 1'b1;
			partial_clause[0][43] 	= 1'b1;
			partial_clause[0][44] 	= ~x[40];
			partial_clause[0][45] 	= 1'b1;
			partial_clause[0][46] 	= 1'b1;
			partial_clause[0][47] 	= 1'b1;
			partial_clause[0][48] 	= 1'b1;
			partial_clause[0][49] 	= 1'b1;
			partial_clause[0][50] 	= 1'b1;
			partial_clause[0][51] 	= 1'b1;
			partial_clause[0][52] 	= ~x[39] & ~x[58];
			partial_clause[0][53] 	= ~x[24];
			partial_clause[0][54] 	= ~x[10];
			partial_clause[0][55] 	= ~x[62];
			partial_clause[0][56] 	= ~x[20] & ~x[24] & ~x[35];
			partial_clause[0][57] 	= ~x[35];
			partial_clause[0][58] 	= 1'b1;
			partial_clause[0][59] 	= ~x[62];
			partial_clause[0][60] 	= ~x[34];
			partial_clause[0][61] 	= ~x[34];
			partial_clause[0][62] 	= 1'b1;
			partial_clause[0][63] 	= 1'b1;
			partial_clause[0][64] 	= ~x[20] & ~x[25] & ~x[44];
			partial_clause[0][65] 	= 1'b1;
			partial_clause[0][66] 	= ~x[37] & ~x[59];
			partial_clause[0][67] 	= ~x[39] & ~x[59];
			partial_clause[0][68] 	= 1'b1;
			partial_clause[0][69] 	= ~x[59];
			partial_clause[0][70] 	= 1'b1;
			partial_clause[0][71] 	= ~x[25] & ~x[36] & ~x[49];
			partial_clause[0][72] 	= ~x[4];
			partial_clause[0][73] 	= ~x[38] & ~x[53];
			partial_clause[0][74] 	= ~x[63];
			partial_clause[0][75] 	= 1'b1;
			partial_clause[0][76] 	= ~x[39];
			partial_clause[0][77] 	= 1'b1;
			partial_clause[0][78] 	= 1'b1;
			partial_clause[0][79] 	= 1'b1;
			partial_clause[0][80] 	= ~x[32];
			partial_clause[0][81] 	= ~x[25];
			partial_clause[0][82] 	= 1'b1;
			partial_clause[0][83] 	= 1'b1;
			partial_clause[0][84] 	= ~x[26] & ~x[47];
			partial_clause[0][85] 	= ~x[24] & ~x[55] & ~x[58];
			partial_clause[0][86] 	= ~x[0] & ~x[44];
			partial_clause[0][87] 	= ~x[4];
			partial_clause[0][88] 	= 1'b1;
			partial_clause[0][89] 	= ~x[45] & ~x[50] & ~x[59];
			partial_clause[0][90] 	= ~x[48] & ~x[59];
			partial_clause[0][91] 	= ~x[18];
			partial_clause[0][92] 	= 1'b1;
			partial_clause[0][93] 	= ~x[50] & ~x[51] & ~x[59];
			partial_clause[0][94] 	= 1'b1;
			partial_clause[0][95] 	= ~x[4] & ~x[34];
			partial_clause[0][96] 	= ~x[48];
			partial_clause[0][97] 	= 1'b1;
			partial_clause[0][98] 	= ~x[9] & ~x[27];
			partial_clause[0][99] 	= ~x[4];
			// Class 1
			partial_clause[1][0] 	= 1'b1;
			partial_clause[1][1] 	= 1'b1;
			partial_clause[1][2] 	= 1'b1;
			partial_clause[1][3] 	= 1'b1;
			partial_clause[1][4] 	= 1'b1;
			partial_clause[1][5] 	= 1'b1;
			partial_clause[1][6] 	= 1'b1;
			partial_clause[1][7] 	= 1'b1;
			partial_clause[1][8] 	= 1'b1;
			partial_clause[1][9] 	= 1'b1;
			partial_clause[1][10] 	= 1'b1;
			partial_clause[1][11] 	= 1'b1;
			partial_clause[1][12] 	= 1'b1;
			partial_clause[1][13] 	= 1'b1;
			partial_clause[1][14] 	= 1'b1;
			partial_clause[1][15] 	= 1'b1;
			partial_clause[1][16] 	= 1'b1;
			partial_clause[1][17] 	= 1'b1;
			partial_clause[1][18] 	= 1'b1;
			partial_clause[1][19] 	= 1'b1;
			partial_clause[1][20] 	= 1'b1;
			partial_clause[1][21] 	= 1'b1;
			partial_clause[1][22] 	= 1'b1;
			partial_clause[1][23] 	= ~x[16];
			partial_clause[1][24] 	= ~x[49];
			partial_clause[1][25] 	= 1'b1;
			partial_clause[1][26] 	= 1'b1;
			partial_clause[1][27] 	= 1'b1;
			partial_clause[1][28] 	= 1'b1;
			partial_clause[1][29] 	= 1'b1;
			partial_clause[1][30] 	= 1'b1;
			partial_clause[1][31] 	= 1'b1;
			partial_clause[1][32] 	= 1'b1;
			partial_clause[1][33] 	= 1'b1;
			partial_clause[1][34] 	= 1'b1;
			partial_clause[1][35] 	= ~x[43];
			partial_clause[1][36] 	= 1'b1;
			partial_clause[1][37] 	= 1'b1;
			partial_clause[1][38] 	= 1'b1;
			partial_clause[1][39] 	= 1'b1;
			partial_clause[1][40] 	= 1'b1;
			partial_clause[1][41] 	= ~x[3];
			partial_clause[1][42] 	= 1'b1;
			partial_clause[1][43] 	= 1'b1;
			partial_clause[1][44] 	= 1'b1;
			partial_clause[1][45] 	= 1'b1;
			partial_clause[1][46] 	= 1'b1;
			partial_clause[1][47] 	= 1'b1;
			partial_clause[1][48] 	= 1'b1;
			partial_clause[1][49] 	= 1'b1;
			partial_clause[1][50] 	= ~x[3] & ~x[36];
			partial_clause[1][51] 	= ~x[60];
			partial_clause[1][52] 	= 1'b1;
			partial_clause[1][53] 	= ~x[32];
			partial_clause[1][54] 	= ~x[28];
			partial_clause[1][55] 	= 1'b1;
			partial_clause[1][56] 	= ~x[20] & ~x[29];
			partial_clause[1][57] 	= ~x[29] & ~x[46];
			partial_clause[1][58] 	= ~x[58];
			partial_clause[1][59] 	= ~x[4] & ~x[11];
			partial_clause[1][60] 	= ~x[25];
			partial_clause[1][61] 	= 1'b1;
			partial_clause[1][62] 	= ~x[26];
			partial_clause[1][63] 	= ~x[36];
			partial_clause[1][64] 	= ~x[4] & ~x[38];
			partial_clause[1][65] 	= ~x[29];
			partial_clause[1][66] 	= ~x[28] & ~x[37];
			partial_clause[1][67] 	= 1'b1;
			partial_clause[1][68] 	= ~x[17];
			partial_clause[1][69] 	= ~x[14];
			partial_clause[1][70] 	= 1'b1;
			partial_clause[1][71] 	= ~x[9];
			partial_clause[1][72] 	= ~x[25] & ~x[53];
			partial_clause[1][73] 	= ~x[18] & ~x[22] & ~x[32];
			partial_clause[1][74] 	= 1'b1;
			partial_clause[1][75] 	= ~x[47];
			partial_clause[1][76] 	= ~x[30];
			partial_clause[1][77] 	= ~x[36] & ~x[43];
			partial_clause[1][78] 	= ~x[0] & ~x[36] & ~x[39];
			partial_clause[1][79] 	= ~x[51] & ~x[55];
			partial_clause[1][80] 	= ~x[18];
			partial_clause[1][81] 	= 1'b1;
			partial_clause[1][82] 	= ~x[9] & ~x[12] & ~x[34];
			partial_clause[1][83] 	= ~x[27] & ~x[51] & ~x[59];
			partial_clause[1][84] 	= 1'b1;
			partial_clause[1][85] 	= ~x[7];
			partial_clause[1][86] 	= ~x[33];
			partial_clause[1][87] 	= ~x[37];
			partial_clause[1][88] 	= ~x[62];
			partial_clause[1][89] 	= ~x[61];
			partial_clause[1][90] 	= ~x[0] & ~x[24] & ~x[55];
			partial_clause[1][91] 	= ~x[16];
			partial_clause[1][92] 	= ~x[32] & ~x[51];
			partial_clause[1][93] 	= ~x[16] & ~x[55];
			partial_clause[1][94] 	= ~x[24];
			partial_clause[1][95] 	= ~x[18] & ~x[35] & ~x[60];
			partial_clause[1][96] 	= ~x[31] & ~x[54];
			partial_clause[1][97] 	= 1'b1;
			partial_clause[1][98] 	= 1'b1;
			partial_clause[1][99] 	= ~x[3] & ~x[25] & ~x[42];
			// Class 2
			partial_clause[2][0] 	= ~x[33];
			partial_clause[2][1] 	= 1'b1;
			partial_clause[2][2] 	= 1'b1;
			partial_clause[2][3] 	= 1'b1;
			partial_clause[2][4] 	= 1'b1;
			partial_clause[2][5] 	= 1'b1;
			partial_clause[2][6] 	= ~x[18] & ~x[25];
			partial_clause[2][7] 	= 1'b1;
			partial_clause[2][8] 	= 1'b1;
			partial_clause[2][9] 	= 1'b1;
			partial_clause[2][10] 	= 1'b1;
			partial_clause[2][11] 	= ~x[46];
			partial_clause[2][12] 	= ~x[14] & ~x[62];
			partial_clause[2][13] 	= 1'b1;
			partial_clause[2][14] 	= 1'b1;
			partial_clause[2][15] 	= 1'b1;
			partial_clause[2][16] 	= ~x[58];
			partial_clause[2][17] 	= 1'b1;
			partial_clause[2][18] 	= ~x[62];
			partial_clause[2][19] 	= 1'b1;
			partial_clause[2][20] 	= 1'b1;
			partial_clause[2][21] 	= 1'b1;
			partial_clause[2][22] 	= 1'b1;
			partial_clause[2][23] 	= ~x[36];
			partial_clause[2][24] 	= 1'b1;
			partial_clause[2][25] 	= 1'b1;
			partial_clause[2][26] 	= ~x[39];
			partial_clause[2][27] 	= 1'b1;
			partial_clause[2][28] 	= 1'b1;
			partial_clause[2][29] 	= 1'b1;
			partial_clause[2][30] 	= ~x[1];
			partial_clause[2][31] 	= 1'b1;
			partial_clause[2][32] 	= ~x[38];
			partial_clause[2][33] 	= 1'b1;
			partial_clause[2][34] 	= 1'b1;
			partial_clause[2][35] 	= ~x[51];
			partial_clause[2][36] 	= 1'b1;
			partial_clause[2][37] 	= ~x[57];
			partial_clause[2][38] 	= 1'b1;
			partial_clause[2][39] 	= 1'b1;
			partial_clause[2][40] 	= ~x[34];
			partial_clause[2][41] 	= 1'b1;
			partial_clause[2][42] 	= 1'b1;
			partial_clause[2][43] 	= 1'b1;
			partial_clause[2][44] 	= 1'b1;
			partial_clause[2][45] 	= 1'b1;
			partial_clause[2][46] 	= ~x[61];
			partial_clause[2][47] 	= 1'b1;
			partial_clause[2][48] 	= 1'b1;
			partial_clause[2][49] 	= 1'b1;
			partial_clause[2][50] 	= 1'b1;
			partial_clause[2][51] 	= 1'b1;
			partial_clause[2][52] 	= 1'b1;
			partial_clause[2][53] 	= 1'b1;
			partial_clause[2][54] 	= 1'b1;
			partial_clause[2][55] 	= 1'b1;
			partial_clause[2][56] 	= ~x[49];
			partial_clause[2][57] 	= 1'b1;
			partial_clause[2][58] 	= ~x[26] & ~x[58];
			partial_clause[2][59] 	= 1'b1;
			partial_clause[2][60] 	= 1'b1;
			partial_clause[2][61] 	= 1'b1;
			partial_clause[2][62] 	= ~x[43];
			partial_clause[2][63] 	= 1'b1;
			partial_clause[2][64] 	= 1'b1;
			partial_clause[2][65] 	= 1'b1;
			partial_clause[2][66] 	= 1'b1;
			partial_clause[2][67] 	= 1'b1;
			partial_clause[2][68] 	= ~x[20];
			partial_clause[2][69] 	= ~x[0];
			partial_clause[2][70] 	= 1'b1;
			partial_clause[2][71] 	= ~x[15] & ~x[33];
			partial_clause[2][72] 	= 1'b1;
			partial_clause[2][73] 	= 1'b1;
			partial_clause[2][74] 	= 1'b1;
			partial_clause[2][75] 	= ~x[22];
			partial_clause[2][76] 	= ~x[9];
			partial_clause[2][77] 	= ~x[43];
			partial_clause[2][78] 	= 1'b1;
			partial_clause[2][79] 	= ~x[46];
			partial_clause[2][80] 	= ~x[26] & ~x[32];
			partial_clause[2][81] 	= ~x[21];
			partial_clause[2][82] 	= 1'b1;
			partial_clause[2][83] 	= 1'b1;
			partial_clause[2][84] 	= 1'b1;
			partial_clause[2][85] 	= 1'b1;
			partial_clause[2][86] 	= 1'b1;
			partial_clause[2][87] 	= 1'b1;
			partial_clause[2][88] 	= ~x[33];
			partial_clause[2][89] 	= 1'b1;
			partial_clause[2][90] 	= ~x[47];
			partial_clause[2][91] 	= 1'b1;
			partial_clause[2][92] 	= ~x[24];
			partial_clause[2][93] 	= 1'b1;
			partial_clause[2][94] 	= 1'b1;
			partial_clause[2][95] 	= 1'b1;
			partial_clause[2][96] 	= 1'b1;
			partial_clause[2][97] 	= 1'b1;
			partial_clause[2][98] 	= ~x[22] & ~x[24] & ~x[55];
			partial_clause[2][99] 	= 1'b1;
			// Class 3
			partial_clause[3][0] 	= 1'b1;
			partial_clause[3][1] 	= ~x[29];
			partial_clause[3][2] 	= 1'b1;
			partial_clause[3][3] 	= ~x[27];
			partial_clause[3][4] 	= 1'b1;
			partial_clause[3][5] 	= 1'b1;
			partial_clause[3][6] 	= 1'b1;
			partial_clause[3][7] 	= ~x[7];
			partial_clause[3][8] 	= 1'b1;
			partial_clause[3][9] 	= 1'b1;
			partial_clause[3][10] 	= 1'b1;
			partial_clause[3][11] 	= ~x[59];
			partial_clause[3][12] 	= ~x[53];
			partial_clause[3][13] 	= 1'b1;
			partial_clause[3][14] 	= 1'b1;
			partial_clause[3][15] 	= 1'b1;
			partial_clause[3][16] 	= 1'b1;
			partial_clause[3][17] 	= 1'b1;
			partial_clause[3][18] 	= ~x[48];
			partial_clause[3][19] 	= 1'b1;
			partial_clause[3][20] 	= 1'b1;
			partial_clause[3][21] 	= 1'b1;
			partial_clause[3][22] 	= ~x[54];
			partial_clause[3][23] 	= 1'b1;
			partial_clause[3][24] 	= 1'b1;
			partial_clause[3][25] 	= 1'b1;
			partial_clause[3][26] 	= 1'b1;
			partial_clause[3][27] 	= ~x[19];
			partial_clause[3][28] 	= ~x[16];
			partial_clause[3][29] 	= 1'b1;
			partial_clause[3][30] 	= 1'b1;
			partial_clause[3][31] 	= 1'b1;
			partial_clause[3][32] 	= ~x[32];
			partial_clause[3][33] 	= 1'b1;
			partial_clause[3][34] 	= 1'b1;
			partial_clause[3][35] 	= ~x[24] & ~x[25];
			partial_clause[3][36] 	= ~x[31];
			partial_clause[3][37] 	= ~x[19];
			partial_clause[3][38] 	= ~x[1];
			partial_clause[3][39] 	= 1'b1;
			partial_clause[3][40] 	= ~x[2] & ~x[25];
			partial_clause[3][41] 	= 1'b1;
			partial_clause[3][42] 	= ~x[50];
			partial_clause[3][43] 	= 1'b1;
			partial_clause[3][44] 	= 1'b1;
			partial_clause[3][45] 	= 1'b1;
			partial_clause[3][46] 	= 1'b1;
			partial_clause[3][47] 	= 1'b1;
			partial_clause[3][48] 	= ~x[27];
			partial_clause[3][49] 	= ~x[16] & ~x[33] & ~x[45];
			partial_clause[3][50] 	= 1'b1;
			partial_clause[3][51] 	= ~x[28];
			partial_clause[3][52] 	= ~x[24] & ~x[31];
			partial_clause[3][53] 	= ~x[10];
			partial_clause[3][54] 	= 1'b1;
			partial_clause[3][55] 	= ~x[9];
			partial_clause[3][56] 	= 1'b1;
			partial_clause[3][57] 	= 1'b1;
			partial_clause[3][58] 	= ~x[18] & ~x[19] & ~x[55];
			partial_clause[3][59] 	= ~x[3] & ~x[45];
			partial_clause[3][60] 	= 1'b1;
			partial_clause[3][61] 	= ~x[11] & ~x[51];
			partial_clause[3][62] 	= 1'b1;
			partial_clause[3][63] 	= ~x[52];
			partial_clause[3][64] 	= 1'b1;
			partial_clause[3][65] 	= 1'b1;
			partial_clause[3][66] 	= ~x[31] & ~x[49];
			partial_clause[3][67] 	= ~x[9] & ~x[37];
			partial_clause[3][68] 	= ~x[5] & ~x[19];
			partial_clause[3][69] 	= 1'b1;
			partial_clause[3][70] 	= ~x[15];
			partial_clause[3][71] 	= 1'b1;
			partial_clause[3][72] 	= ~x[9] & ~x[30];
			partial_clause[3][73] 	= ~x[48];
			partial_clause[3][74] 	= ~x[12] & ~x[20] & ~x[31];
			partial_clause[3][75] 	= 1'b1;
			partial_clause[3][76] 	= 1'b1;
			partial_clause[3][77] 	= ~x[33];
			partial_clause[3][78] 	= ~x[25] & ~x[44];
			partial_clause[3][79] 	= 1'b1;
			partial_clause[3][80] 	= ~x[40];
			partial_clause[3][81] 	= ~x[28] & ~x[33] & ~x[41];
			partial_clause[3][82] 	= ~x[15] & ~x[22];
			partial_clause[3][83] 	= 1'b1;
			partial_clause[3][84] 	= 1'b1;
			partial_clause[3][85] 	= ~x[45];
			partial_clause[3][86] 	= ~x[4];
			partial_clause[3][87] 	= ~x[60];
			partial_clause[3][88] 	= ~x[4];
			partial_clause[3][89] 	= 1'b1;
			partial_clause[3][90] 	= ~x[23];
			partial_clause[3][91] 	= ~x[34];
			partial_clause[3][92] 	= ~x[44];
			partial_clause[3][93] 	= 1'b1;
			partial_clause[3][94] 	= ~x[30] & ~x[56];
			partial_clause[3][95] 	= ~x[16] & ~x[34] & ~x[43] & ~x[61];
			partial_clause[3][96] 	= 1'b1;
			partial_clause[3][97] 	= 1'b1;
			partial_clause[3][98] 	= ~x[31];
			partial_clause[3][99] 	= ~x[11] & ~x[34];
			// Class 4
			partial_clause[4][0] 	= 1'b1;
			partial_clause[4][1] 	= ~x[34];
			partial_clause[4][2] 	= ~x[43];
			partial_clause[4][3] 	= 1'b1;
			partial_clause[4][4] 	= ~x[6];
			partial_clause[4][5] 	= 1'b1;
			partial_clause[4][6] 	= 1'b1;
			partial_clause[4][7] 	= 1'b1;
			partial_clause[4][8] 	= ~x[55];
			partial_clause[4][9] 	= 1'b1;
			partial_clause[4][10] 	= 1'b1;
			partial_clause[4][11] 	= 1'b1;
			partial_clause[4][12] 	= 1'b1;
			partial_clause[4][13] 	= ~x[22];
			partial_clause[4][14] 	= 1'b1;
			partial_clause[4][15] 	= 1'b1;
			partial_clause[4][16] 	= 1'b1;
			partial_clause[4][17] 	= 1'b1;
			partial_clause[4][18] 	= 1'b1;
			partial_clause[4][19] 	= 1'b1;
			partial_clause[4][20] 	= 1'b1;
			partial_clause[4][21] 	= ~x[30];
			partial_clause[4][22] 	= ~x[56];
			partial_clause[4][23] 	= ~x[28];
			partial_clause[4][24] 	= 1'b1;
			partial_clause[4][25] 	= 1'b1;
			partial_clause[4][26] 	= ~x[43];
			partial_clause[4][27] 	= 1'b1;
			partial_clause[4][28] 	= 1'b1;
			partial_clause[4][29] 	= ~x[29];
			partial_clause[4][30] 	= 1'b1;
			partial_clause[4][31] 	= ~x[1] & ~x[11];
			partial_clause[4][32] 	= 1'b1;
			partial_clause[4][33] 	= 1'b1;
			partial_clause[4][34] 	= 1'b1;
			partial_clause[4][35] 	= 1'b1;
			partial_clause[4][36] 	= ~x[6] & ~x[63];
			partial_clause[4][37] 	= 1'b1;
			partial_clause[4][38] 	= 1'b1;
			partial_clause[4][39] 	= 1'b1;
			partial_clause[4][40] 	= 1'b1;
			partial_clause[4][41] 	= 1'b1;
			partial_clause[4][42] 	= ~x[31];
			partial_clause[4][43] 	= 1'b1;
			partial_clause[4][44] 	= 1'b1;
			partial_clause[4][45] 	= 1'b1;
			partial_clause[4][46] 	= 1'b1;
			partial_clause[4][47] 	= ~x[38];
			partial_clause[4][48] 	= 1'b1;
			partial_clause[4][49] 	= 1'b1;
			partial_clause[4][50] 	= ~x[6];
			partial_clause[4][51] 	= 1'b1;
			partial_clause[4][52] 	= 1'b1;
			partial_clause[4][53] 	= ~x[36] & ~x[43] & ~x[49];
			partial_clause[4][54] 	= 1'b1;
			partial_clause[4][55] 	= 1'b1;
			partial_clause[4][56] 	= ~x[14] & ~x[23];
			partial_clause[4][57] 	= ~x[4] & ~x[52];
			partial_clause[4][58] 	= ~x[31] & ~x[62];
			partial_clause[4][59] 	= 1'b1;
			partial_clause[4][60] 	= 1'b1;
			partial_clause[4][61] 	= ~x[43];
			partial_clause[4][62] 	= 1'b1;
			partial_clause[4][63] 	= ~x[15] & ~x[56];
			partial_clause[4][64] 	= ~x[43];
			partial_clause[4][65] 	= ~x[18] & ~x[27];
			partial_clause[4][66] 	= ~x[20] & ~x[46] & ~x[50] & ~x[58];
			partial_clause[4][67] 	= 1'b1;
			partial_clause[4][68] 	= ~x[58];
			partial_clause[4][69] 	= ~x[27] & ~x[55];
			partial_clause[4][70] 	= ~x[0] & ~x[15] & ~x[58] & ~x[63];
			partial_clause[4][71] 	= 1'b1;
			partial_clause[4][72] 	= ~x[18] & ~x[24];
			partial_clause[4][73] 	= 1'b1;
			partial_clause[4][74] 	= ~x[12] & ~x[49];
			partial_clause[4][75] 	= ~x[33] & ~x[56];
			partial_clause[4][76] 	= 1'b1;
			partial_clause[4][77] 	= ~x[27];
			partial_clause[4][78] 	= ~x[62];
			partial_clause[4][79] 	= ~x[44];
			partial_clause[4][80] 	= ~x[9] & ~x[14];
			partial_clause[4][81] 	= ~x[2];
			partial_clause[4][82] 	= ~x[2] & ~x[16] & ~x[34];
			partial_clause[4][83] 	= 1'b1;
			partial_clause[4][84] 	= 1'b1;
			partial_clause[4][85] 	= ~x[0];
			partial_clause[4][86] 	= 1'b1;
			partial_clause[4][87] 	= ~x[15];
			partial_clause[4][88] 	= ~x[8] & ~x[11] & ~x[54] & ~x[55];
			partial_clause[4][89] 	= ~x[37] & ~x[42] & ~x[57];
			partial_clause[4][90] 	= ~x[7] & ~x[41];
			partial_clause[4][91] 	= ~x[3] & ~x[5];
			partial_clause[4][92] 	= ~x[27] & ~x[33];
			partial_clause[4][93] 	= ~x[14];
			partial_clause[4][94] 	= ~x[6];
			partial_clause[4][95] 	= ~x[53];
			partial_clause[4][96] 	= 1'b1;
			partial_clause[4][97] 	= 1'b1;
			partial_clause[4][98] 	= ~x[16] & ~x[52];
			partial_clause[4][99] 	= ~x[31];
			// Class 5
			partial_clause[5][0] 	= 1'b1;
			partial_clause[5][1] 	= ~x[22] & ~x[60];
			partial_clause[5][2] 	= 1'b1;
			partial_clause[5][3] 	= 1'b1;
			partial_clause[5][4] 	= 1'b1;
			partial_clause[5][5] 	= ~x[45];
			partial_clause[5][6] 	= 1'b1;
			partial_clause[5][7] 	= ~x[41];
			partial_clause[5][8] 	= 1'b1;
			partial_clause[5][9] 	= 1'b1;
			partial_clause[5][10] 	= 1'b1;
			partial_clause[5][11] 	= 1'b1;
			partial_clause[5][12] 	= 1'b1;
			partial_clause[5][13] 	= 1'b1;
			partial_clause[5][14] 	= 1'b1;
			partial_clause[5][15] 	= 1'b1;
			partial_clause[5][16] 	= 1'b1;
			partial_clause[5][17] 	= ~x[9] & ~x[57];
			partial_clause[5][18] 	= 1'b1;
			partial_clause[5][19] 	= ~x[36];
			partial_clause[5][20] 	= 1'b1;
			partial_clause[5][21] 	= 1'b1;
			partial_clause[5][22] 	= 1'b1;
			partial_clause[5][23] 	= 1'b1;
			partial_clause[5][24] 	= 1'b1;
			partial_clause[5][25] 	= 1'b1;
			partial_clause[5][26] 	= 1'b1;
			partial_clause[5][27] 	= 1'b1;
			partial_clause[5][28] 	= 1'b1;
			partial_clause[5][29] 	= 1'b1;
			partial_clause[5][30] 	= ~x[35] & ~x[49];
			partial_clause[5][31] 	= 1'b1;
			partial_clause[5][32] 	= 1'b1;
			partial_clause[5][33] 	= 1'b1;
			partial_clause[5][34] 	= ~x[37];
			partial_clause[5][35] 	= 1'b1;
			partial_clause[5][36] 	= ~x[5];
			partial_clause[5][37] 	= 1'b1;
			partial_clause[5][38] 	= 1'b1;
			partial_clause[5][39] 	= 1'b1;
			partial_clause[5][40] 	= 1'b1;
			partial_clause[5][41] 	= 1'b1;
			partial_clause[5][42] 	= 1'b1;
			partial_clause[5][43] 	= ~x[56];
			partial_clause[5][44] 	= 1'b1;
			partial_clause[5][45] 	= 1'b1;
			partial_clause[5][46] 	= 1'b1;
			partial_clause[5][47] 	= 1'b1;
			partial_clause[5][48] 	= 1'b1;
			partial_clause[5][49] 	= 1'b1;
			partial_clause[5][50] 	= 1'b1;
			partial_clause[5][51] 	= 1'b1;
			partial_clause[5][52] 	= ~x[12] & ~x[58];
			partial_clause[5][53] 	= ~x[19];
			partial_clause[5][54] 	= ~x[12];
			partial_clause[5][55] 	= ~x[20] & ~x[42];
			partial_clause[5][56] 	= ~x[34];
			partial_clause[5][57] 	= ~x[39];
			partial_clause[5][58] 	= ~x[18] & ~x[44];
			partial_clause[5][59] 	= 1'b1;
			partial_clause[5][60] 	= 1'b1;
			partial_clause[5][61] 	= ~x[46];
			partial_clause[5][62] 	= 1'b1;
			partial_clause[5][63] 	= ~x[62];
			partial_clause[5][64] 	= ~x[22];
			partial_clause[5][65] 	= ~x[40];
			partial_clause[5][66] 	= ~x[41];
			partial_clause[5][67] 	= 1'b1;
			partial_clause[5][68] 	= 1'b1;
			partial_clause[5][69] 	= 1'b1;
			partial_clause[5][70] 	= ~x[3];
			partial_clause[5][71] 	= 1'b1;
			partial_clause[5][72] 	= 1'b1;
			partial_clause[5][73] 	= 1'b1;
			partial_clause[5][74] 	= 1'b1;
			partial_clause[5][75] 	= ~x[23];
			partial_clause[5][76] 	= 1'b1;
			partial_clause[5][77] 	= 1'b1;
			partial_clause[5][78] 	= ~x[15] & ~x[19];
			partial_clause[5][79] 	= 1'b1;
			partial_clause[5][80] 	= 1'b1;
			partial_clause[5][81] 	= 1'b1;
			partial_clause[5][82] 	= ~x[7];
			partial_clause[5][83] 	= 1'b1;
			partial_clause[5][84] 	= 1'b1;
			partial_clause[5][85] 	= ~x[53];
			partial_clause[5][86] 	= ~x[31];
			partial_clause[5][87] 	= ~x[13];
			partial_clause[5][88] 	= ~x[25];
			partial_clause[5][89] 	= 1'b1;
			partial_clause[5][90] 	= 1'b1;
			partial_clause[5][91] 	= ~x[44];
			partial_clause[5][92] 	= 1'b1;
			partial_clause[5][93] 	= 1'b1;
			partial_clause[5][94] 	= ~x[6];
			partial_clause[5][95] 	= ~x[23] & ~x[55];
			partial_clause[5][96] 	= 1'b1;
			partial_clause[5][97] 	= 1'b1;
			partial_clause[5][98] 	= 1'b1;
			partial_clause[5][99] 	= ~x[23];
			// Class 6
			partial_clause[6][0] 	= 1'b1;
			partial_clause[6][1] 	= 1'b1;
			partial_clause[6][2] 	= 1'b1;
			partial_clause[6][3] 	= 1'b1;
			partial_clause[6][4] 	= 1'b1;
			partial_clause[6][5] 	= 1'b1;
			partial_clause[6][6] 	= ~x[34];
			partial_clause[6][7] 	= ~x[12];
			partial_clause[6][8] 	= 1'b1;
			partial_clause[6][9] 	= ~x[33];
			partial_clause[6][10] 	= 1'b1;
			partial_clause[6][11] 	= 1'b1;
			partial_clause[6][12] 	= 1'b1;
			partial_clause[6][13] 	= ~x[18];
			partial_clause[6][14] 	= 1'b1;
			partial_clause[6][15] 	= 1'b1;
			partial_clause[6][16] 	= ~x[52];
			partial_clause[6][17] 	= 1'b1;
			partial_clause[6][18] 	= 1'b1;
			partial_clause[6][19] 	= ~x[13];
			partial_clause[6][20] 	= 1'b1;
			partial_clause[6][21] 	= 1'b1;
			partial_clause[6][22] 	= 1'b1;
			partial_clause[6][23] 	= 1'b1;
			partial_clause[6][24] 	= 1'b1;
			partial_clause[6][25] 	= 1'b1;
			partial_clause[6][26] 	= ~x[28];
			partial_clause[6][27] 	= 1'b1;
			partial_clause[6][28] 	= 1'b1;
			partial_clause[6][29] 	= 1'b1;
			partial_clause[6][30] 	= 1'b1;
			partial_clause[6][31] 	= ~x[14];
			partial_clause[6][32] 	= 1'b1;
			partial_clause[6][33] 	= 1'b1;
			partial_clause[6][34] 	= ~x[28];
			partial_clause[6][35] 	= ~x[12];
			partial_clause[6][36] 	= 1'b1;
			partial_clause[6][37] 	= 1'b1;
			partial_clause[6][38] 	= 1'b1;
			partial_clause[6][39] 	= ~x[47];
			partial_clause[6][40] 	= 1'b1;
			partial_clause[6][41] 	= 1'b1;
			partial_clause[6][42] 	= 1'b1;
			partial_clause[6][43] 	= 1'b1;
			partial_clause[6][44] 	= 1'b1;
			partial_clause[6][45] 	= ~x[37];
			partial_clause[6][46] 	= ~x[52];
			partial_clause[6][47] 	= 1'b1;
			partial_clause[6][48] 	= ~x[38];
			partial_clause[6][49] 	= 1'b1;
			partial_clause[6][50] 	= 1'b1;
			partial_clause[6][51] 	= ~x[48];
			partial_clause[6][52] 	= ~x[0] & ~x[17];
			partial_clause[6][53] 	= ~x[35];
			partial_clause[6][54] 	= 1'b1;
			partial_clause[6][55] 	= 1'b1;
			partial_clause[6][56] 	= 1'b1;
			partial_clause[6][57] 	= 1'b1;
			partial_clause[6][58] 	= ~x[5];
			partial_clause[6][59] 	= ~x[33];
			partial_clause[6][60] 	= ~x[62];
			partial_clause[6][61] 	= 1'b1;
			partial_clause[6][62] 	= 1'b1;
			partial_clause[6][63] 	= ~x[49] & ~x[50];
			partial_clause[6][64] 	= 1'b1;
			partial_clause[6][65] 	= ~x[2];
			partial_clause[6][66] 	= 1'b1;
			partial_clause[6][67] 	= 1'b1;
			partial_clause[6][68] 	= 1'b1;
			partial_clause[6][69] 	= ~x[36];
			partial_clause[6][70] 	= ~x[24];
			partial_clause[6][71] 	= ~x[25];
			partial_clause[6][72] 	= 1'b1;
			partial_clause[6][73] 	= ~x[18] & ~x[49];
			partial_clause[6][74] 	= ~x[49];
			partial_clause[6][75] 	= ~x[10] & ~x[43];
			partial_clause[6][76] 	= 1'b1;
			partial_clause[6][77] 	= 1'b1;
			partial_clause[6][78] 	= ~x[50];
			partial_clause[6][79] 	= 1'b1;
			partial_clause[6][80] 	= 1'b1;
			partial_clause[6][81] 	= 1'b1;
			partial_clause[6][82] 	= ~x[57];
			partial_clause[6][83] 	= ~x[5];
			partial_clause[6][84] 	= 1'b1;
			partial_clause[6][85] 	= 1'b1;
			partial_clause[6][86] 	= ~x[13];
			partial_clause[6][87] 	= ~x[34];
			partial_clause[6][88] 	= ~x[9] & ~x[38];
			partial_clause[6][89] 	= 1'b1;
			partial_clause[6][90] 	= ~x[40];
			partial_clause[6][91] 	= ~x[11];
			partial_clause[6][92] 	= ~x[24] & ~x[49];
			partial_clause[6][93] 	= 1'b1;
			partial_clause[6][94] 	= ~x[47];
			partial_clause[6][95] 	= 1'b1;
			partial_clause[6][96] 	= 1'b1;
			partial_clause[6][97] 	= 1'b1;
			partial_clause[6][98] 	= ~x[38];
			partial_clause[6][99] 	= 1'b1;
			// Class 7
			partial_clause[7][0] 	= 1'b1;
			partial_clause[7][1] 	= 1'b1;
			partial_clause[7][2] 	= 1'b1;
			partial_clause[7][3] 	= 1'b1;
			partial_clause[7][4] 	= ~x[20];
			partial_clause[7][5] 	= 1'b1;
			partial_clause[7][6] 	= 1'b1;
			partial_clause[7][7] 	= 1'b1;
			partial_clause[7][8] 	= 1'b1;
			partial_clause[7][9] 	= 1'b1;
			partial_clause[7][10] 	= 1'b1;
			partial_clause[7][11] 	= 1'b1;
			partial_clause[7][12] 	= ~x[47];
			partial_clause[7][13] 	= ~x[33];
			partial_clause[7][14] 	= 1'b1;
			partial_clause[7][15] 	= 1'b1;
			partial_clause[7][16] 	= 1'b1;
			partial_clause[7][17] 	= ~x[4];
			partial_clause[7][18] 	= 1'b1;
			partial_clause[7][19] 	= 1'b1;
			partial_clause[7][20] 	= 1'b1;
			partial_clause[7][21] 	= 1'b1;
			partial_clause[7][22] 	= 1'b1;
			partial_clause[7][23] 	= 1'b1;
			partial_clause[7][24] 	= 1'b1;
			partial_clause[7][25] 	= 1'b1;
			partial_clause[7][26] 	= 1'b1;
			partial_clause[7][27] 	= 1'b1;
			partial_clause[7][28] 	= 1'b1;
			partial_clause[7][29] 	= 1'b1;
			partial_clause[7][30] 	= 1'b1;
			partial_clause[7][31] 	= 1'b1;
			partial_clause[7][32] 	= 1'b1;
			partial_clause[7][33] 	= ~x[34];
			partial_clause[7][34] 	= 1'b1;
			partial_clause[7][35] 	= 1'b1;
			partial_clause[7][36] 	= 1'b1;
			partial_clause[7][37] 	= 1'b1;
			partial_clause[7][38] 	= 1'b1;
			partial_clause[7][39] 	= ~x[12];
			partial_clause[7][40] 	= 1'b1;
			partial_clause[7][41] 	= ~x[47];
			partial_clause[7][42] 	= 1'b1;
			partial_clause[7][43] 	= 1'b1;
			partial_clause[7][44] 	= 1'b1;
			partial_clause[7][45] 	= ~x[0];
			partial_clause[7][46] 	= 1'b1;
			partial_clause[7][47] 	= ~x[56];
			partial_clause[7][48] 	= ~x[9];
			partial_clause[7][49] 	= 1'b1;
			partial_clause[7][50] 	= 1'b1;
			partial_clause[7][51] 	= 1'b1;
			partial_clause[7][52] 	= ~x[10];
			partial_clause[7][53] 	= ~x[6] & ~x[59];
			partial_clause[7][54] 	= 1'b1;
			partial_clause[7][55] 	= 1'b1;
			partial_clause[7][56] 	= ~x[34];
			partial_clause[7][57] 	= 1'b1;
			partial_clause[7][58] 	= ~x[56];
			partial_clause[7][59] 	= 1'b1;
			partial_clause[7][60] 	= ~x[26];
			partial_clause[7][61] 	= 1'b1;
			partial_clause[7][62] 	= ~x[46];
			partial_clause[7][63] 	= 1'b1;
			partial_clause[7][64] 	= 1'b1;
			partial_clause[7][65] 	= ~x[3] & ~x[32];
			partial_clause[7][66] 	= 1'b1;
			partial_clause[7][67] 	= 1'b1;
			partial_clause[7][68] 	= ~x[18] & ~x[62];
			partial_clause[7][69] 	= 1'b1;
			partial_clause[7][70] 	= ~x[40];
			partial_clause[7][71] 	= ~x[37];
			partial_clause[7][72] 	= 1'b1;
			partial_clause[7][73] 	= 1'b1;
			partial_clause[7][74] 	= 1'b1;
			partial_clause[7][75] 	= 1'b1;
			partial_clause[7][76] 	= 1'b1;
			partial_clause[7][77] 	= 1'b1;
			partial_clause[7][78] 	= 1'b1;
			partial_clause[7][79] 	= ~x[2] & ~x[24];
			partial_clause[7][80] 	= ~x[2];
			partial_clause[7][81] 	= 1'b1;
			partial_clause[7][82] 	= 1'b1;
			partial_clause[7][83] 	= 1'b1;
			partial_clause[7][84] 	= 1'b1;
			partial_clause[7][85] 	= 1'b1;
			partial_clause[7][86] 	= ~x[19] & ~x[40];
			partial_clause[7][87] 	= 1'b1;
			partial_clause[7][88] 	= 1'b1;
			partial_clause[7][89] 	= 1'b1;
			partial_clause[7][90] 	= ~x[60];
			partial_clause[7][91] 	= 1'b1;
			partial_clause[7][92] 	= 1'b1;
			partial_clause[7][93] 	= 1'b1;
			partial_clause[7][94] 	= ~x[19];
			partial_clause[7][95] 	= ~x[60];
			partial_clause[7][96] 	= 1'b1;
			partial_clause[7][97] 	= 1'b1;
			partial_clause[7][98] 	= 1'b1;
			partial_clause[7][99] 	= 1'b1;
			// Class 8
			partial_clause[8][0] 	= ~x[4] & ~x[58];
			partial_clause[8][1] 	= 1'b1;
			partial_clause[8][2] 	= 1'b1;
			partial_clause[8][3] 	= 1'b1;
			partial_clause[8][4] 	= 1'b1;
			partial_clause[8][5] 	= 1'b1;
			partial_clause[8][6] 	= ~x[19] & ~x[37];
			partial_clause[8][7] 	= 1'b1;
			partial_clause[8][8] 	= 1'b1;
			partial_clause[8][9] 	= ~x[33];
			partial_clause[8][10] 	= 1'b1;
			partial_clause[8][11] 	= ~x[56];
			partial_clause[8][12] 	= ~x[13];
			partial_clause[8][13] 	= ~x[14] & ~x[38];
			partial_clause[8][14] 	= ~x[26];
			partial_clause[8][15] 	= ~x[14];
			partial_clause[8][16] 	= 1'b1;
			partial_clause[8][17] 	= ~x[35] & ~x[55];
			partial_clause[8][18] 	= 1'b1;
			partial_clause[8][19] 	= ~x[40];
			partial_clause[8][20] 	= 1'b1;
			partial_clause[8][21] 	= 1'b1;
			partial_clause[8][22] 	= ~x[47];
			partial_clause[8][23] 	= ~x[18];
			partial_clause[8][24] 	= 1'b1;
			partial_clause[8][25] 	= ~x[54];
			partial_clause[8][26] 	= 1'b1;
			partial_clause[8][27] 	= 1'b1;
			partial_clause[8][28] 	= ~x[43];
			partial_clause[8][29] 	= ~x[23];
			partial_clause[8][30] 	= ~x[49];
			partial_clause[8][31] 	= 1'b1;
			partial_clause[8][32] 	= ~x[32];
			partial_clause[8][33] 	= ~x[8] & ~x[42];
			partial_clause[8][34] 	= 1'b1;
			partial_clause[8][35] 	= ~x[48];
			partial_clause[8][36] 	= ~x[21];
			partial_clause[8][37] 	= 1'b1;
			partial_clause[8][38] 	= 1'b1;
			partial_clause[8][39] 	= 1'b1;
			partial_clause[8][40] 	= 1'b1;
			partial_clause[8][41] 	= 1'b1;
			partial_clause[8][42] 	= 1'b1;
			partial_clause[8][43] 	= 1'b1;
			partial_clause[8][44] 	= 1'b1;
			partial_clause[8][45] 	= 1'b1;
			partial_clause[8][46] 	= 1'b1;
			partial_clause[8][47] 	= 1'b1;
			partial_clause[8][48] 	= ~x[21];
			partial_clause[8][49] 	= 1'b1;
			partial_clause[8][50] 	= ~x[36] & ~x[37];
			partial_clause[8][51] 	= ~x[60];
			partial_clause[8][52] 	= ~x[43];
			partial_clause[8][53] 	= ~x[15];
			partial_clause[8][54] 	= ~x[17];
			partial_clause[8][55] 	= ~x[38] & ~x[60];
			partial_clause[8][56] 	= 1'b1;
			partial_clause[8][57] 	= ~x[38];
			partial_clause[8][58] 	= ~x[39];
			partial_clause[8][59] 	= ~x[3] & ~x[4] & ~x[20];
			partial_clause[8][60] 	= 1'b1;
			partial_clause[8][61] 	= 1'b1;
			partial_clause[8][62] 	= ~x[10] & ~x[23];
			partial_clause[8][63] 	= ~x[50];
			partial_clause[8][64] 	= ~x[37];
			partial_clause[8][65] 	= ~x[9] & ~x[10] & ~x[56];
			partial_clause[8][66] 	= ~x[27];
			partial_clause[8][67] 	= ~x[12];
			partial_clause[8][68] 	= ~x[61];
			partial_clause[8][69] 	= ~x[5];
			partial_clause[8][70] 	= ~x[41];
			partial_clause[8][71] 	= ~x[0] & ~x[24];
			partial_clause[8][72] 	= ~x[11];
			partial_clause[8][73] 	= 1'b1;
			partial_clause[8][74] 	= ~x[7] & ~x[33];
			partial_clause[8][75] 	= 1'b1;
			partial_clause[8][76] 	= 1'b1;
			partial_clause[8][77] 	= 1'b1;
			partial_clause[8][78] 	= ~x[44];
			partial_clause[8][79] 	= 1'b1;
			partial_clause[8][80] 	= ~x[32];
			partial_clause[8][81] 	= 1'b1;
			partial_clause[8][82] 	= ~x[11] & ~x[48] & ~x[57];
			partial_clause[8][83] 	= 1'b1;
			partial_clause[8][84] 	= ~x[2];
			partial_clause[8][85] 	= ~x[6];
			partial_clause[8][86] 	= 1'b1;
			partial_clause[8][87] 	= 1'b1;
			partial_clause[8][88] 	= 1'b1;
			partial_clause[8][89] 	= 1'b1;
			partial_clause[8][90] 	= ~x[23] & ~x[45];
			partial_clause[8][91] 	= ~x[30] & ~x[46];
			partial_clause[8][92] 	= ~x[53];
			partial_clause[8][93] 	= ~x[34];
			partial_clause[8][94] 	= ~x[25];
			partial_clause[8][95] 	= ~x[29];
			partial_clause[8][96] 	= ~x[1] & ~x[60];
			partial_clause[8][97] 	= ~x[2];
			partial_clause[8][98] 	= ~x[49];
			partial_clause[8][99] 	= 1'b1;
			// Class 9
			partial_clause[9][0] 	= 1'b1;
			partial_clause[9][1] 	= 1'b1;
			partial_clause[9][2] 	= 1'b1;
			partial_clause[9][3] 	= 1'b1;
			partial_clause[9][4] 	= 1'b1;
			partial_clause[9][5] 	= 1'b1;
			partial_clause[9][6] 	= 1'b1;
			partial_clause[9][7] 	= 1'b1;
			partial_clause[9][8] 	= 1'b1;
			partial_clause[9][9] 	= 1'b1;
			partial_clause[9][10] 	= 1'b1;
			partial_clause[9][11] 	= 1'b1;
			partial_clause[9][12] 	= 1'b1;
			partial_clause[9][13] 	= ~x[54];
			partial_clause[9][14] 	= 1'b1;
			partial_clause[9][15] 	= 1'b1;
			partial_clause[9][16] 	= 1'b1;
			partial_clause[9][17] 	= 1'b1;
			partial_clause[9][18] 	= 1'b1;
			partial_clause[9][19] 	= 1'b1;
			partial_clause[9][20] 	= ~x[9] & ~x[52];
			partial_clause[9][21] 	= 1'b1;
			partial_clause[9][22] 	= 1'b1;
			partial_clause[9][23] 	= 1'b1;
			partial_clause[9][24] 	= 1'b1;
			partial_clause[9][25] 	= ~x[0];
			partial_clause[9][26] 	= 1'b1;
			partial_clause[9][27] 	= 1'b1;
			partial_clause[9][28] 	= 1'b1;
			partial_clause[9][29] 	= 1'b1;
			partial_clause[9][30] 	= 1'b1;
			partial_clause[9][31] 	= 1'b1;
			partial_clause[9][32] 	= 1'b1;
			partial_clause[9][33] 	= 1'b1;
			partial_clause[9][34] 	= 1'b1;
			partial_clause[9][35] 	= 1'b1;
			partial_clause[9][36] 	= ~x[14];
			partial_clause[9][37] 	= ~x[21];
			partial_clause[9][38] 	= 1'b1;
			partial_clause[9][39] 	= 1'b1;
			partial_clause[9][40] 	= 1'b1;
			partial_clause[9][41] 	= ~x[2];
			partial_clause[9][42] 	= 1'b1;
			partial_clause[9][43] 	= ~x[5];
			partial_clause[9][44] 	= 1'b1;
			partial_clause[9][45] 	= ~x[24];
			partial_clause[9][46] 	= 1'b1;
			partial_clause[9][47] 	= 1'b1;
			partial_clause[9][48] 	= 1'b1;
			partial_clause[9][49] 	= ~x[62];
			partial_clause[9][50] 	= 1'b1;
			partial_clause[9][51] 	= 1'b1;
			partial_clause[9][52] 	= ~x[35];
			partial_clause[9][53] 	= 1'b1;
			partial_clause[9][54] 	= ~x[15] & ~x[55];
			partial_clause[9][55] 	= 1'b1;
			partial_clause[9][56] 	= 1'b1;
			partial_clause[9][57] 	= ~x[16] & ~x[58];
			partial_clause[9][58] 	= ~x[1];
			partial_clause[9][59] 	= ~x[62];
			partial_clause[9][60] 	= ~x[35];
			partial_clause[9][61] 	= 1'b1;
			partial_clause[9][62] 	= 1'b1;
			partial_clause[9][63] 	= 1'b1;
			partial_clause[9][64] 	= 1'b1;
			partial_clause[9][65] 	= 1'b1;
			partial_clause[9][66] 	= 1'b1;
			partial_clause[9][67] 	= 1'b1;
			partial_clause[9][68] 	= 1'b1;
			partial_clause[9][69] 	= 1'b1;
			partial_clause[9][70] 	= 1'b1;
			partial_clause[9][71] 	= 1'b1;
			partial_clause[9][72] 	= ~x[26];
			partial_clause[9][73] 	= ~x[26];
			partial_clause[9][74] 	= ~x[45];
			partial_clause[9][75] 	= 1'b1;
			partial_clause[9][76] 	= ~x[22];
			partial_clause[9][77] 	= 1'b1;
			partial_clause[9][78] 	= 1'b1;
			partial_clause[9][79] 	= ~x[4];
			partial_clause[9][80] 	= 1'b1;
			partial_clause[9][81] 	= 1'b1;
			partial_clause[9][82] 	= ~x[35] & ~x[37];
			partial_clause[9][83] 	= ~x[51];
			partial_clause[9][84] 	= ~x[15];
			partial_clause[9][85] 	= 1'b1;
			partial_clause[9][86] 	= ~x[18];
			partial_clause[9][87] 	= ~x[51];
			partial_clause[9][88] 	= ~x[21];
			partial_clause[9][89] 	= 1'b1;
			partial_clause[9][90] 	= ~x[52];
			partial_clause[9][91] 	= 1'b1;
			partial_clause[9][92] 	= ~x[6] & ~x[11];
			partial_clause[9][93] 	= 1'b1;
			partial_clause[9][94] 	= 1'b1;
			partial_clause[9][95] 	= 1'b1;
			partial_clause[9][96] 	= 1'b1;
			partial_clause[9][97] 	= 1'b1;
			partial_clause[9][98] 	= ~x[24];
			partial_clause[9][99] 	= ~x[55];
		end
	end
endmodule


module HCB_1 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & ~x[5];
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & ~x[53];
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & ~x[32];
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & ~x[9];
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & ~x[13];
			partial_clause[0][20] 	= partial_clause_prev[0][20] & ~x[55];
			partial_clause[0][21] 	= partial_clause_prev[0][21] & ~x[12] & ~x[32];
			partial_clause[0][22] 	= partial_clause_prev[0][22] & ~x[47];
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & ~x[44];
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & ~x[16];
			partial_clause[0][32] 	= partial_clause_prev[0][32] & ~x[32];
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & ~x[7];
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & ~x[18];
			partial_clause[0][40] 	= partial_clause_prev[0][40] & ~x[21] & ~x[26];
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & ~x[15] & ~x[57];
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & ~x[31];
			partial_clause[0][50] 	= partial_clause_prev[0][50] & ~x[25] & ~x[44];
			partial_clause[0][51] 	= partial_clause_prev[0][51] & ~x[22];
			partial_clause[0][52] 	= partial_clause_prev[0][52] & ~x[18];
			partial_clause[0][53] 	= partial_clause_prev[0][53] & ~x[13];
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & ~x[51];
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & ~x[2];
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & ~x[49];
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & ~x[17] & ~x[51];
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & ~x[1];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & ~x[47];
			partial_clause[0][74] 	= partial_clause_prev[0][74] & ~x[43] & ~x[52];
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & ~x[19];
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & ~x[51];
			partial_clause[0][79] 	= partial_clause_prev[0][79] & ~x[17];
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & ~x[40];
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & ~x[25];
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & ~x[18] & ~x[26];
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & ~x[18] & ~x[51];
			partial_clause[0][94] 	= partial_clause_prev[0][94] & ~x[28];
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & ~x[27];
			partial_clause[0][97] 	= partial_clause_prev[0][97] & ~x[23];
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & ~x[50];
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & ~x[35];
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & ~x[11];
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & ~x[28];
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & ~x[55];
			partial_clause[1][29] 	= partial_clause_prev[1][29] & ~x[3];
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & ~x[55];
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & ~x[7];
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & ~x[28];
			partial_clause[1][52] 	= partial_clause_prev[1][52] & ~x[52];
			partial_clause[1][53] 	= partial_clause_prev[1][53] & ~x[13] & ~x[46];
			partial_clause[1][54] 	= partial_clause_prev[1][54] & ~x[26] & ~x[52];
			partial_clause[1][55] 	= partial_clause_prev[1][55] & ~x[22] & ~x[50];
			partial_clause[1][56] 	= partial_clause_prev[1][56] & ~x[26];
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & ~x[51];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & ~x[18];
			partial_clause[1][61] 	= partial_clause_prev[1][61] & ~x[2] & ~x[45];
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & ~x[11];
			partial_clause[1][64] 	= partial_clause_prev[1][64] & ~x[24];
			partial_clause[1][65] 	= partial_clause_prev[1][65] & ~x[20];
			partial_clause[1][66] 	= partial_clause_prev[1][66] & ~x[27];
			partial_clause[1][67] 	= partial_clause_prev[1][67] & ~x[24] & ~x[46];
			partial_clause[1][68] 	= partial_clause_prev[1][68] & ~x[2];
			partial_clause[1][69] 	= partial_clause_prev[1][69] & ~x[45];
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & ~x[16] & ~x[18] & ~x[58] & ~x[59];
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & ~x[20];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & ~x[26] & ~x[48];
			partial_clause[1][76] 	= partial_clause_prev[1][76] & ~x[18];
			partial_clause[1][77] 	= partial_clause_prev[1][77] & ~x[25];
			partial_clause[1][78] 	= partial_clause_prev[1][78] & ~x[41];
			partial_clause[1][79] 	= partial_clause_prev[1][79] & ~x[16] & ~x[51];
			partial_clause[1][80] 	= partial_clause_prev[1][80] & ~x[27] & ~x[55];
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & ~x[9];
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & ~x[45] & ~x[47] & ~x[49];
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & ~x[21] & ~x[25];
			partial_clause[1][89] 	= partial_clause_prev[1][89] & ~x[7] & ~x[49];
			partial_clause[1][90] 	= partial_clause_prev[1][90] & ~x[19];
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & ~x[1];
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & ~x[17];
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & ~x[23] & ~x[51];
			partial_clause[1][98] 	= partial_clause_prev[1][98] & ~x[12];
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & ~x[47];
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & ~x[50];
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & ~x[40];
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & ~x[49];
			partial_clause[2][18] 	= partial_clause_prev[2][18] & ~x[46];
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & ~x[44];
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & ~x[21] & ~x[44];
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & ~x[16];
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & ~x[12];
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & ~x[48];
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & ~x[52];
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & ~x[47];
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & ~x[59];
			partial_clause[2][52] 	= partial_clause_prev[2][52] & ~x[56] & ~x[59];
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & ~x[60];
			partial_clause[2][55] 	= partial_clause_prev[2][55] & ~x[31] & ~x[32];
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & ~x[36] & ~x[60];
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & ~x[56] & ~x[58];
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & ~x[58];
			partial_clause[2][63] 	= partial_clause_prev[2][63] & ~x[63];
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & 1'b1;
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & ~x[57];
			partial_clause[2][68] 	= partial_clause_prev[2][68] & ~x[25] & ~x[28];
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & ~x[60];
			partial_clause[2][73] 	= partial_clause_prev[2][73] & ~x[31] & ~x[32] & ~x[58];
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & ~x[31] & ~x[60];
			partial_clause[2][76] 	= partial_clause_prev[2][76] & ~x[33];
			partial_clause[2][77] 	= partial_clause_prev[2][77] & ~x[3] & ~x[20] & ~x[59];
			partial_clause[2][78] 	= partial_clause_prev[2][78] & ~x[62] & ~x[63];
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & ~x[61];
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & ~x[57];
			partial_clause[2][85] 	= partial_clause_prev[2][85] & ~x[61] & ~x[62];
			partial_clause[2][86] 	= partial_clause_prev[2][86] & ~x[29];
			partial_clause[2][87] 	= partial_clause_prev[2][87] & ~x[60] & ~x[61];
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & ~x[4] & ~x[58];
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & ~x[61];
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & ~x[57] & ~x[60];
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & ~x[16];
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & ~x[22];
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & ~x[18];
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & ~x[42];
			partial_clause[3][7] 	= partial_clause_prev[3][7] & ~x[8];
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & ~x[18];
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & ~x[18];
			partial_clause[3][18] 	= partial_clause_prev[3][18] & ~x[13];
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & ~x[36];
			partial_clause[3][25] 	= partial_clause_prev[3][25] & ~x[16];
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & ~x[16] & ~x[18] & ~x[40];
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & ~x[46];
			partial_clause[3][34] 	= partial_clause_prev[3][34] & ~x[1];
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & ~x[28];
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & ~x[56];
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & ~x[18];
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & ~x[54];
			partial_clause[3][63] 	= partial_clause_prev[3][63] & ~x[60];
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & 1'b1;
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & ~x[48];
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & ~x[48] & ~x[56];
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & ~x[22] & ~x[28] & ~x[31] & ~x[59];
			partial_clause[3][76] 	= partial_clause_prev[3][76] & ~x[23];
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & ~x[60];
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & ~x[49];
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & ~x[60];
			partial_clause[3][88] 	= partial_clause_prev[3][88] & ~x[28];
			partial_clause[3][89] 	= partial_clause_prev[3][89] & ~x[26];
			partial_clause[3][90] 	= partial_clause_prev[3][90] & ~x[49];
			partial_clause[3][91] 	= partial_clause_prev[3][91] & ~x[16] & ~x[19];
			partial_clause[3][92] 	= partial_clause_prev[3][92] & ~x[16];
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & ~x[46] & ~x[50];
			partial_clause[3][98] 	= partial_clause_prev[3][98] & ~x[33];
			partial_clause[3][99] 	= partial_clause_prev[3][99] & ~x[60];
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & ~x[3] & ~x[58];
			partial_clause[4][1] 	= partial_clause_prev[4][1] & ~x[30] & ~x[33];
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & ~x[32] & ~x[62] & ~x[63];
			partial_clause[4][4] 	= partial_clause_prev[4][4] & ~x[23] & ~x[63];
			partial_clause[4][5] 	= partial_clause_prev[4][5] & ~x[36] & ~x[62];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & ~x[3] & ~x[33] & ~x[40];
			partial_clause[4][7] 	= partial_clause_prev[4][7] & ~x[17] & ~x[62];
			partial_clause[4][8] 	= partial_clause_prev[4][8] & ~x[49];
			partial_clause[4][9] 	= partial_clause_prev[4][9] & ~x[33] & ~x[53] & ~x[62];
			partial_clause[4][10] 	= partial_clause_prev[4][10] & ~x[34] & ~x[60] & ~x[63];
			partial_clause[4][11] 	= partial_clause_prev[4][11] & ~x[32] & ~x[57] & ~x[63];
			partial_clause[4][12] 	= partial_clause_prev[4][12] & ~x[62];
			partial_clause[4][13] 	= partial_clause_prev[4][13] & ~x[31] & ~x[32];
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & ~x[62];
			partial_clause[4][16] 	= partial_clause_prev[4][16] & ~x[3];
			partial_clause[4][17] 	= partial_clause_prev[4][17] & ~x[58] & ~x[60] & ~x[63];
			partial_clause[4][18] 	= partial_clause_prev[4][18] & ~x[33] & ~x[53];
			partial_clause[4][19] 	= partial_clause_prev[4][19] & ~x[24] & ~x[61];
			partial_clause[4][20] 	= partial_clause_prev[4][20] & ~x[33] & ~x[34];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & ~x[63];
			partial_clause[4][22] 	= partial_clause_prev[4][22] & ~x[6] & ~x[59];
			partial_clause[4][23] 	= partial_clause_prev[4][23] & ~x[62];
			partial_clause[4][24] 	= partial_clause_prev[4][24] & ~x[5] & ~x[6] & ~x[63];
			partial_clause[4][25] 	= partial_clause_prev[4][25] & ~x[32] & ~x[35] & ~x[61];
			partial_clause[4][26] 	= partial_clause_prev[4][26] & ~x[34] & ~x[63];
			partial_clause[4][27] 	= partial_clause_prev[4][27] & ~x[33] & ~x[50];
			partial_clause[4][28] 	= partial_clause_prev[4][28] & ~x[9] & ~x[35] & ~x[37] & ~x[60] & ~x[63];
			partial_clause[4][29] 	= partial_clause_prev[4][29] & ~x[33] & ~x[35];
			partial_clause[4][30] 	= partial_clause_prev[4][30] & ~x[32] & ~x[38] & ~x[61];
			partial_clause[4][31] 	= partial_clause_prev[4][31] & ~x[61];
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[33];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & ~x[31] & ~x[62];
			partial_clause[4][34] 	= partial_clause_prev[4][34] & ~x[59];
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & ~x[63];
			partial_clause[4][37] 	= partial_clause_prev[4][37] & ~x[29] & ~x[60];
			partial_clause[4][38] 	= partial_clause_prev[4][38] & ~x[33] & ~x[34];
			partial_clause[4][39] 	= partial_clause_prev[4][39] & ~x[59] & ~x[62];
			partial_clause[4][40] 	= partial_clause_prev[4][40] & ~x[6] & ~x[21] & ~x[32] & ~x[63];
			partial_clause[4][41] 	= partial_clause_prev[4][41] & ~x[34] & ~x[62];
			partial_clause[4][42] 	= partial_clause_prev[4][42] & ~x[34] & ~x[60] & ~x[63];
			partial_clause[4][43] 	= partial_clause_prev[4][43] & ~x[5] & ~x[31] & ~x[52];
			partial_clause[4][44] 	= partial_clause_prev[4][44] & ~x[13];
			partial_clause[4][45] 	= partial_clause_prev[4][45] & ~x[33];
			partial_clause[4][46] 	= partial_clause_prev[4][46] & ~x[36];
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & ~x[34] & ~x[45] & ~x[59];
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[35] & ~x[37];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & ~x[11] & ~x[16];
			partial_clause[4][52] 	= partial_clause_prev[4][52] & ~x[24] & ~x[54];
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & ~x[0];
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & ~x[51];
			partial_clause[4][59] 	= partial_clause_prev[4][59] & ~x[18];
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & ~x[8];
			partial_clause[4][63] 	= partial_clause_prev[4][63] & ~x[13];
			partial_clause[4][64] 	= partial_clause_prev[4][64] & ~x[15];
			partial_clause[4][65] 	= partial_clause_prev[4][65] & ~x[18];
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & ~x[19];
			partial_clause[4][68] 	= partial_clause_prev[4][68] & ~x[52];
			partial_clause[4][69] 	= partial_clause_prev[4][69] & ~x[29];
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & ~x[49];
			partial_clause[4][75] 	= partial_clause_prev[4][75] & ~x[20];
			partial_clause[4][76] 	= partial_clause_prev[4][76] & ~x[24];
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & ~x[4];
			partial_clause[4][79] 	= partial_clause_prev[4][79] & ~x[28];
			partial_clause[4][80] 	= partial_clause_prev[4][80] & ~x[1] & ~x[25];
			partial_clause[4][81] 	= partial_clause_prev[4][81] & ~x[46] & ~x[53];
			partial_clause[4][82] 	= partial_clause_prev[4][82] & ~x[16];
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & ~x[0];
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & ~x[6] & ~x[14] & ~x[15];
			partial_clause[4][90] 	= partial_clause_prev[4][90] & ~x[12] & ~x[26] & ~x[52];
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & ~x[16];
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & ~x[6] & ~x[46];
			partial_clause[4][98] 	= partial_clause_prev[4][98] & ~x[22];
			partial_clause[4][99] 	= partial_clause_prev[4][99] & ~x[3] & ~x[4];
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & ~x[61] & ~x[63];
			partial_clause[5][1] 	= partial_clause_prev[5][1] & ~x[34];
			partial_clause[5][2] 	= partial_clause_prev[5][2] & ~x[40] & ~x[51] & ~x[63];
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & ~x[40];
			partial_clause[5][5] 	= partial_clause_prev[5][5] & ~x[20] & ~x[34] & ~x[49];
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & ~x[8];
			partial_clause[5][9] 	= partial_clause_prev[5][9] & ~x[41] & ~x[55];
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & ~x[36];
			partial_clause[5][12] 	= partial_clause_prev[5][12] & ~x[33];
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & ~x[61];
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & ~x[55];
			partial_clause[5][19] 	= partial_clause_prev[5][19] & ~x[35];
			partial_clause[5][20] 	= partial_clause_prev[5][20] & ~x[58];
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & ~x[37] & ~x[49];
			partial_clause[5][23] 	= partial_clause_prev[5][23] & ~x[9];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & ~x[10];
			partial_clause[5][26] 	= partial_clause_prev[5][26] & ~x[7];
			partial_clause[5][27] 	= partial_clause_prev[5][27] & ~x[6];
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & ~x[9] & ~x[17];
			partial_clause[5][33] 	= partial_clause_prev[5][33] & ~x[55];
			partial_clause[5][34] 	= partial_clause_prev[5][34] & ~x[36];
			partial_clause[5][35] 	= partial_clause_prev[5][35] & ~x[34];
			partial_clause[5][36] 	= partial_clause_prev[5][36] & ~x[33] & ~x[34];
			partial_clause[5][37] 	= partial_clause_prev[5][37] & ~x[38];
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & ~x[19];
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & ~x[30];
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & ~x[36];
			partial_clause[5][45] 	= partial_clause_prev[5][45] & ~x[8] & ~x[39] & ~x[55];
			partial_clause[5][46] 	= partial_clause_prev[5][46] & ~x[38];
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & ~x[39];
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & ~x[24];
			partial_clause[5][61] 	= partial_clause_prev[5][61] & ~x[27];
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & ~x[42];
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & ~x[49];
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & ~x[16];
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & ~x[2];
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & ~x[2];
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & ~x[23] & ~x[25];
			partial_clause[5][78] 	= partial_clause_prev[5][78] & ~x[51];
			partial_clause[5][79] 	= partial_clause_prev[5][79] & ~x[27];
			partial_clause[5][80] 	= partial_clause_prev[5][80] & ~x[1];
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & ~x[15];
			partial_clause[5][83] 	= partial_clause_prev[5][83] & ~x[23];
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & ~x[18];
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & ~x[42];
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & ~x[10];
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & ~x[41] & ~x[51];
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & ~x[22] & ~x[27];
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & ~x[21];
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & ~x[2] & ~x[28] & ~x[29] & ~x[30] & ~x[35] & ~x[37];
			partial_clause[6][51] 	= partial_clause_prev[6][51] & ~x[31] & ~x[34] & ~x[36] & ~x[38] & ~x[39] & ~x[40];
			partial_clause[6][52] 	= partial_clause_prev[6][52] & ~x[28] & ~x[43];
			partial_clause[6][53] 	= partial_clause_prev[6][53] & ~x[6] & ~x[9] & ~x[30];
			partial_clause[6][54] 	= partial_clause_prev[6][54] & ~x[0] & ~x[4] & ~x[25] & ~x[34] & ~x[35] & ~x[36] & ~x[38];
			partial_clause[6][55] 	= partial_clause_prev[6][55] & ~x[35] & ~x[38] & ~x[40];
			partial_clause[6][56] 	= partial_clause_prev[6][56] & ~x[12] & ~x[32] & ~x[34] & ~x[36] & ~x[38];
			partial_clause[6][57] 	= partial_clause_prev[6][57] & ~x[33] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[58];
			partial_clause[6][58] 	= partial_clause_prev[6][58] & ~x[30] & ~x[32] & ~x[35] & ~x[36] & ~x[37] & ~x[39] & ~x[42];
			partial_clause[6][59] 	= partial_clause_prev[6][59] & ~x[3] & ~x[40] & ~x[44];
			partial_clause[6][60] 	= partial_clause_prev[6][60] & ~x[36] & ~x[39] & ~x[50];
			partial_clause[6][61] 	= partial_clause_prev[6][61] & ~x[30] & ~x[35] & ~x[52] & ~x[55];
			partial_clause[6][62] 	= partial_clause_prev[6][62] & ~x[9] & ~x[31] & ~x[35] & ~x[39];
			partial_clause[6][63] 	= partial_clause_prev[6][63] & ~x[3] & ~x[34] & ~x[35] & ~x[37] & ~x[38];
			partial_clause[6][64] 	= partial_clause_prev[6][64] & ~x[33] & ~x[38] & ~x[40] & ~x[41];
			partial_clause[6][65] 	= partial_clause_prev[6][65] & ~x[30] & ~x[33] & ~x[36] & ~x[37] & ~x[39] & ~x[57];
			partial_clause[6][66] 	= partial_clause_prev[6][66] & ~x[35] & ~x[43] & ~x[49] & ~x[51];
			partial_clause[6][67] 	= partial_clause_prev[6][67] & ~x[16] & ~x[35] & ~x[37] & ~x[38] & ~x[40] & ~x[44];
			partial_clause[6][68] 	= partial_clause_prev[6][68] & ~x[32] & ~x[33] & ~x[36] & ~x[40] & ~x[57];
			partial_clause[6][69] 	= partial_clause_prev[6][69] & ~x[0] & ~x[31] & ~x[32] & ~x[34] & ~x[35] & ~x[39] & ~x[40];
			partial_clause[6][70] 	= partial_clause_prev[6][70] & ~x[0];
			partial_clause[6][71] 	= partial_clause_prev[6][71] & ~x[10] & ~x[40];
			partial_clause[6][72] 	= partial_clause_prev[6][72] & ~x[2] & ~x[33] & ~x[34] & ~x[36] & ~x[38];
			partial_clause[6][73] 	= partial_clause_prev[6][73] & ~x[2] & ~x[28] & ~x[32] & ~x[37] & ~x[38] & ~x[40];
			partial_clause[6][74] 	= partial_clause_prev[6][74] & ~x[3] & ~x[35] & ~x[40];
			partial_clause[6][75] 	= partial_clause_prev[6][75] & ~x[28] & ~x[29] & ~x[34];
			partial_clause[6][76] 	= partial_clause_prev[6][76] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[41];
			partial_clause[6][77] 	= partial_clause_prev[6][77] & ~x[31] & ~x[34] & ~x[35] & ~x[37] & ~x[39];
			partial_clause[6][78] 	= partial_clause_prev[6][78] & ~x[37];
			partial_clause[6][79] 	= partial_clause_prev[6][79] & ~x[33] & ~x[36] & ~x[38] & ~x[58];
			partial_clause[6][80] 	= partial_clause_prev[6][80] & ~x[35] & ~x[37] & ~x[39] & ~x[40] & ~x[43];
			partial_clause[6][81] 	= partial_clause_prev[6][81] & ~x[4] & ~x[10] & ~x[27] & ~x[30] & ~x[32] & ~x[35] & ~x[37] & ~x[39];
			partial_clause[6][82] 	= partial_clause_prev[6][82] & ~x[31] & ~x[38];
			partial_clause[6][83] 	= partial_clause_prev[6][83] & ~x[17];
			partial_clause[6][84] 	= partial_clause_prev[6][84] & ~x[29] & ~x[30] & ~x[33] & ~x[38];
			partial_clause[6][85] 	= partial_clause_prev[6][85] & ~x[6] & ~x[32] & ~x[33] & ~x[36] & ~x[37];
			partial_clause[6][86] 	= partial_clause_prev[6][86] & ~x[5] & ~x[33] & ~x[35] & ~x[37];
			partial_clause[6][87] 	= partial_clause_prev[6][87] & ~x[40] & ~x[42];
			partial_clause[6][88] 	= partial_clause_prev[6][88] & ~x[3] & ~x[33] & ~x[35] & ~x[36] & ~x[37] & ~x[39];
			partial_clause[6][89] 	= partial_clause_prev[6][89] & ~x[9] & ~x[12] & ~x[35] & ~x[37];
			partial_clause[6][90] 	= partial_clause_prev[6][90] & ~x[55] & ~x[57];
			partial_clause[6][91] 	= partial_clause_prev[6][91] & ~x[14] & ~x[33];
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & ~x[3] & ~x[4] & ~x[33] & ~x[35] & ~x[36] & ~x[38] & ~x[39] & ~x[41];
			partial_clause[6][94] 	= partial_clause_prev[6][94] & ~x[5] & ~x[36] & ~x[37] & ~x[38];
			partial_clause[6][95] 	= partial_clause_prev[6][95] & ~x[5] & ~x[34] & ~x[36] & ~x[38];
			partial_clause[6][96] 	= partial_clause_prev[6][96] & ~x[2] & ~x[32] & ~x[35] & ~x[36] & ~x[37] & ~x[40];
			partial_clause[6][97] 	= partial_clause_prev[6][97] & ~x[31] & ~x[33] & ~x[35] & ~x[36] & ~x[37] & ~x[38];
			partial_clause[6][98] 	= partial_clause_prev[6][98] & ~x[38] & ~x[40];
			partial_clause[6][99] 	= partial_clause_prev[6][99] & ~x[31] & ~x[36] & ~x[38] & ~x[39];
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & ~x[31];
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & ~x[15];
			partial_clause[7][3] 	= partial_clause_prev[7][3] & ~x[57];
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & ~x[61];
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & ~x[63];
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & ~x[36];
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & ~x[62];
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & ~x[60];
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & ~x[59];
			partial_clause[7][25] 	= partial_clause_prev[7][25] & ~x[61];
			partial_clause[7][26] 	= partial_clause_prev[7][26] & ~x[31] & ~x[63];
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & ~x[13];
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & ~x[50];
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & ~x[63];
			partial_clause[7][35] 	= partial_clause_prev[7][35] & ~x[62];
			partial_clause[7][36] 	= partial_clause_prev[7][36] & ~x[57];
			partial_clause[7][37] 	= partial_clause_prev[7][37] & ~x[37];
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & ~x[62];
			partial_clause[7][40] 	= partial_clause_prev[7][40] & ~x[63];
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & ~x[60] & ~x[63];
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & ~x[62];
			partial_clause[7][49] 	= partial_clause_prev[7][49] & ~x[61];
			partial_clause[7][50] 	= partial_clause_prev[7][50] & ~x[53];
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & ~x[9] & ~x[46];
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & ~x[27];
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & ~x[1] & ~x[19] & ~x[25];
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & ~x[0] & ~x[25];
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & ~x[37];
			partial_clause[8][2] 	= partial_clause_prev[8][2] & ~x[39];
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & ~x[34];
			partial_clause[8][6] 	= partial_clause_prev[8][6] & ~x[8];
			partial_clause[8][7] 	= partial_clause_prev[8][7] & ~x[15] & ~x[19] & ~x[27] & ~x[34] & ~x[58];
			partial_clause[8][8] 	= partial_clause_prev[8][8] & ~x[18] & ~x[32];
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & ~x[10];
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & ~x[58];
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & ~x[51];
			partial_clause[8][15] 	= partial_clause_prev[8][15] & ~x[39];
			partial_clause[8][16] 	= partial_clause_prev[8][16] & ~x[35];
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & ~x[21];
			partial_clause[8][19] 	= partial_clause_prev[8][19] & ~x[16] & ~x[29] & ~x[44];
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & ~x[20];
			partial_clause[8][22] 	= partial_clause_prev[8][22] & ~x[6];
			partial_clause[8][23] 	= partial_clause_prev[8][23] & ~x[38];
			partial_clause[8][24] 	= partial_clause_prev[8][24] & ~x[41] & ~x[42] & ~x[59];
			partial_clause[8][25] 	= partial_clause_prev[8][25] & ~x[7];
			partial_clause[8][26] 	= partial_clause_prev[8][26] & ~x[36] & ~x[59];
			partial_clause[8][27] 	= partial_clause_prev[8][27] & ~x[45];
			partial_clause[8][28] 	= partial_clause_prev[8][28] & ~x[36];
			partial_clause[8][29] 	= partial_clause_prev[8][29] & ~x[18] & ~x[37] & ~x[48];
			partial_clause[8][30] 	= partial_clause_prev[8][30] & ~x[36];
			partial_clause[8][31] 	= partial_clause_prev[8][31] & ~x[8] & ~x[26];
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & ~x[16] & ~x[35] & ~x[59];
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & ~x[50];
			partial_clause[8][36] 	= partial_clause_prev[8][36] & ~x[52];
			partial_clause[8][37] 	= partial_clause_prev[8][37] & ~x[59];
			partial_clause[8][38] 	= partial_clause_prev[8][38] & ~x[21] & ~x[28];
			partial_clause[8][39] 	= partial_clause_prev[8][39] & ~x[35];
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & ~x[42];
			partial_clause[8][42] 	= partial_clause_prev[8][42] & ~x[24];
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & ~x[32] & ~x[36];
			partial_clause[8][46] 	= partial_clause_prev[8][46] & ~x[48];
			partial_clause[8][47] 	= partial_clause_prev[8][47] & ~x[7] & ~x[30];
			partial_clause[8][48] 	= partial_clause_prev[8][48] & ~x[33];
			partial_clause[8][49] 	= partial_clause_prev[8][49] & ~x[35];
			partial_clause[8][50] 	= partial_clause_prev[8][50] & ~x[47];
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & ~x[18] & ~x[24];
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & ~x[41];
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & ~x[2];
			partial_clause[8][60] 	= partial_clause_prev[8][60] & ~x[48];
			partial_clause[8][61] 	= partial_clause_prev[8][61] & ~x[44];
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & ~x[13];
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & ~x[52];
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & ~x[24] & ~x[25] & ~x[49];
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & ~x[17];
			partial_clause[8][75] 	= partial_clause_prev[8][75] & ~x[13];
			partial_clause[8][76] 	= partial_clause_prev[8][76] & ~x[48];
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & ~x[10] & ~x[23] & ~x[53];
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & ~x[18];
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & ~x[1];
			partial_clause[8][85] 	= partial_clause_prev[8][85] & ~x[48];
			partial_clause[8][86] 	= partial_clause_prev[8][86] & ~x[52];
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & ~x[2] & ~x[50];
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & ~x[25];
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & ~x[19];
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & ~x[25];
			partial_clause[8][97] 	= partial_clause_prev[8][97] & ~x[52];
			partial_clause[8][98] 	= partial_clause_prev[8][98] & ~x[44];
			partial_clause[8][99] 	= partial_clause_prev[8][99] & ~x[49];
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & ~x[42];
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & ~x[34];
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & ~x[62];
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & ~x[11];
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & ~x[62];
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & ~x[60];
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & ~x[6];
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & 1'b1;
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & ~x[40];
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & ~x[47] & ~x[52];
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & ~x[61];
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & ~x[60];
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & ~x[43] & ~x[48];
			partial_clause[9][53] 	= partial_clause_prev[9][53] & ~x[42];
			partial_clause[9][54] 	= partial_clause_prev[9][54] & ~x[23];
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & ~x[45];
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & ~x[49];
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & ~x[16] & ~x[17];
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & ~x[25];
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & ~x[18];
			partial_clause[9][88] 	= partial_clause_prev[9][88] & ~x[48];
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & ~x[54];
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
		end
	end
endmodule


module HCB_2 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & ~x[40];
			partial_clause[0][6] 	= partial_clause_prev[0][6] & ~x[19];
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & ~x[45];
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & ~x[18];
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & x[56];
			partial_clause[0][16] 	= partial_clause_prev[0][16] & ~x[43];
			partial_clause[0][17] 	= partial_clause_prev[0][17] & ~x[44];
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & ~x[41];
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & ~x[13] & ~x[42];
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & ~x[16];
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & ~x[45];
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & ~x[16];
			partial_clause[0][34] 	= partial_clause_prev[0][34] & ~x[7] & ~x[16] & ~x[46];
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & ~x[46];
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & ~x[10];
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & ~x[8] & ~x[20];
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & ~x[13];
			partial_clause[0][52] 	= partial_clause_prev[0][52] & ~x[14] & ~x[40];
			partial_clause[0][53] 	= partial_clause_prev[0][53] & ~x[12] & ~x[14];
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & ~x[14];
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & ~x[12];
			partial_clause[0][66] 	= partial_clause_prev[0][66] & ~x[14];
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & ~x[16];
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & ~x[17];
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & ~x[10];
			partial_clause[0][83] 	= partial_clause_prev[0][83] & ~x[13];
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & ~x[41];
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & ~x[37];
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & ~x[40];
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & ~x[15];
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[21] & ~x[48];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & ~x[49];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & ~x[49];
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & ~x[22];
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & ~x[49] & ~x[50];
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & ~x[47];
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & ~x[22];
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & ~x[49];
			partial_clause[1][19] 	= partial_clause_prev[1][19] & ~x[22];
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & ~x[21] & ~x[50];
			partial_clause[1][22] 	= partial_clause_prev[1][22] & ~x[50];
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & ~x[13];
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & ~x[49];
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & ~x[36];
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & ~x[47];
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & ~x[48];
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & ~x[49];
			partial_clause[1][48] 	= partial_clause_prev[1][48] & ~x[5] & ~x[61];
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & ~x[18] & ~x[39];
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & ~x[16];
			partial_clause[1][53] 	= partial_clause_prev[1][53] & ~x[7];
			partial_clause[1][54] 	= partial_clause_prev[1][54] & ~x[43];
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & ~x[10];
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & 1'b1;
			partial_clause[1][59] 	= partial_clause_prev[1][59] & ~x[42];
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & ~x[13] & ~x[37];
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & ~x[40];
			partial_clause[1][74] 	= partial_clause_prev[1][74] & 1'b1;
			partial_clause[1][75] 	= partial_clause_prev[1][75] & ~x[40];
			partial_clause[1][76] 	= partial_clause_prev[1][76] & ~x[5] & ~x[9];
			partial_clause[1][77] 	= partial_clause_prev[1][77] & ~x[40];
			partial_clause[1][78] 	= partial_clause_prev[1][78] & ~x[38];
			partial_clause[1][79] 	= partial_clause_prev[1][79] & ~x[37];
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & ~x[8];
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & ~x[4] & ~x[6];
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & ~x[14];
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & ~x[41];
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & x[26];
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & ~x[10];
			partial_clause[2][6] 	= partial_clause_prev[2][6] & ~x[11];
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & ~x[11];
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & x[26];
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & ~x[44];
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & ~x[39];
			partial_clause[2][22] 	= partial_clause_prev[2][22] & ~x[15];
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & ~x[14];
			partial_clause[2][26] 	= partial_clause_prev[2][26] & x[25];
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & x[26];
			partial_clause[2][29] 	= partial_clause_prev[2][29] & x[26];
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & x[25];
			partial_clause[2][32] 	= partial_clause_prev[2][32] & x[25];
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & ~x[40];
			partial_clause[2][37] 	= partial_clause_prev[2][37] & x[26];
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & x[28];
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & x[25];
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & x[26];
			partial_clause[2][44] 	= partial_clause_prev[2][44] & ~x[9];
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & ~x[48];
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & ~x[22] & ~x[23];
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & ~x[24];
			partial_clause[2][60] 	= partial_clause_prev[2][60] & ~x[23];
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & ~x[14];
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & ~x[46];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & ~x[22];
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & ~x[12];
			partial_clause[2][69] 	= partial_clause_prev[2][69] & ~x[17];
			partial_clause[2][70] 	= partial_clause_prev[2][70] & ~x[47];
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & ~x[20] & ~x[21] & ~x[48];
			partial_clause[2][84] 	= partial_clause_prev[2][84] & ~x[20];
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & ~x[37];
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & ~x[49];
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & ~x[23];
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & ~x[23];
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & ~x[5];
			partial_clause[3][1] 	= partial_clause_prev[3][1] & ~x[35];
			partial_clause[3][2] 	= partial_clause_prev[3][2] & ~x[40];
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & ~x[12];
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & x[52];
			partial_clause[3][8] 	= partial_clause_prev[3][8] & ~x[35];
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & ~x[5] & ~x[13];
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & ~x[36];
			partial_clause[3][16] 	= partial_clause_prev[3][16] & ~x[13];
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & x[53];
			partial_clause[3][19] 	= partial_clause_prev[3][19] & ~x[10] & ~x[12] & ~x[63];
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & ~x[63];
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & ~x[63];
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & ~x[35];
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & ~x[7];
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & ~x[63];
			partial_clause[3][37] 	= partial_clause_prev[3][37] & ~x[6];
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & x[55];
			partial_clause[3][43] 	= partial_clause_prev[3][43] & ~x[36];
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & ~x[63];
			partial_clause[3][48] 	= partial_clause_prev[3][48] & ~x[12] & x[55];
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & ~x[44];
			partial_clause[3][51] 	= partial_clause_prev[3][51] & ~x[11] & ~x[25] & ~x[50];
			partial_clause[3][52] 	= partial_clause_prev[3][52] & ~x[14];
			partial_clause[3][53] 	= partial_clause_prev[3][53] & ~x[18];
			partial_clause[3][54] 	= partial_clause_prev[3][54] & ~x[48];
			partial_clause[3][55] 	= partial_clause_prev[3][55] & ~x[45];
			partial_clause[3][56] 	= partial_clause_prev[3][56] & ~x[22] & ~x[48];
			partial_clause[3][57] 	= partial_clause_prev[3][57] & ~x[46];
			partial_clause[3][58] 	= partial_clause_prev[3][58] & ~x[11];
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & ~x[45];
			partial_clause[3][62] 	= partial_clause_prev[3][62] & ~x[12];
			partial_clause[3][63] 	= partial_clause_prev[3][63] & ~x[52] & ~x[53];
			partial_clause[3][64] 	= partial_clause_prev[3][64] & ~x[11] & ~x[22] & ~x[50];
			partial_clause[3][65] 	= partial_clause_prev[3][65] & 1'b1;
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & ~x[17] & ~x[45];
			partial_clause[3][68] 	= partial_clause_prev[3][68] & ~x[22];
			partial_clause[3][69] 	= partial_clause_prev[3][69] & ~x[6];
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & ~x[24] & ~x[52];
			partial_clause[3][72] 	= partial_clause_prev[3][72] & ~x[13];
			partial_clause[3][73] 	= partial_clause_prev[3][73] & ~x[49];
			partial_clause[3][74] 	= partial_clause_prev[3][74] & ~x[41];
			partial_clause[3][75] 	= partial_clause_prev[3][75] & ~x[23];
			partial_clause[3][76] 	= partial_clause_prev[3][76] & ~x[19];
			partial_clause[3][77] 	= partial_clause_prev[3][77] & ~x[12] & ~x[26] & ~x[44] & ~x[54];
			partial_clause[3][78] 	= partial_clause_prev[3][78] & ~x[22];
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & ~x[19] & ~x[22] & ~x[51];
			partial_clause[3][81] 	= partial_clause_prev[3][81] & ~x[20];
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & ~x[24] & ~x[49];
			partial_clause[3][84] 	= partial_clause_prev[3][84] & ~x[13] & ~x[23] & ~x[50];
			partial_clause[3][85] 	= partial_clause_prev[3][85] & ~x[49];
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & ~x[44] & ~x[50];
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & ~x[24];
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & ~x[48];
			partial_clause[3][92] 	= partial_clause_prev[3][92] & ~x[24] & ~x[51];
			partial_clause[3][93] 	= partial_clause_prev[3][93] & ~x[22] & ~x[50];
			partial_clause[3][94] 	= partial_clause_prev[3][94] & ~x[19];
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & ~x[48];
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & ~x[24] & ~x[51];
			partial_clause[3][99] 	= partial_clause_prev[3][99] & ~x[24] & ~x[51];
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & ~x[27] & ~x[54];
			partial_clause[4][1] 	= partial_clause_prev[4][1] & ~x[28];
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & ~x[55];
			partial_clause[4][5] 	= partial_clause_prev[4][5] & ~x[55];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & ~x[27];
			partial_clause[4][7] 	= partial_clause_prev[4][7] & ~x[54];
			partial_clause[4][8] 	= partial_clause_prev[4][8] & ~x[26] & ~x[27];
			partial_clause[4][9] 	= partial_clause_prev[4][9] & ~x[54];
			partial_clause[4][10] 	= partial_clause_prev[4][10] & ~x[55];
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & ~x[54];
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & ~x[16];
			partial_clause[4][15] 	= partial_clause_prev[4][15] & ~x[13] & ~x[54];
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & ~x[27];
			partial_clause[4][18] 	= partial_clause_prev[4][18] & ~x[26] & ~x[54];
			partial_clause[4][19] 	= partial_clause_prev[4][19] & ~x[54];
			partial_clause[4][20] 	= partial_clause_prev[4][20] & ~x[55];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & ~x[55];
			partial_clause[4][25] 	= partial_clause_prev[4][25] & ~x[55];
			partial_clause[4][26] 	= partial_clause_prev[4][26] & ~x[55];
			partial_clause[4][27] 	= partial_clause_prev[4][27] & ~x[26];
			partial_clause[4][28] 	= partial_clause_prev[4][28] & ~x[55];
			partial_clause[4][29] 	= partial_clause_prev[4][29] & ~x[26];
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & ~x[0] & ~x[55];
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[26];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & ~x[55];
			partial_clause[4][34] 	= partial_clause_prev[4][34] & ~x[53];
			partial_clause[4][35] 	= partial_clause_prev[4][35] & ~x[55];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & ~x[55];
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & ~x[27];
			partial_clause[4][39] 	= partial_clause_prev[4][39] & ~x[54];
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & ~x[55];
			partial_clause[4][42] 	= partial_clause_prev[4][42] & ~x[56];
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & ~x[55];
			partial_clause[4][45] 	= partial_clause_prev[4][45] & ~x[27];
			partial_clause[4][46] 	= partial_clause_prev[4][46] & ~x[56];
			partial_clause[4][47] 	= partial_clause_prev[4][47] & ~x[53];
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[27];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & x[54] & x[56];
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & x[53] & x[55];
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & ~x[43];
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & x[54] & x[56];
			partial_clause[4][62] 	= partial_clause_prev[4][62] & x[55];
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & ~x[15] & ~x[62] & ~x[63];
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & x[55];
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & ~x[12] & ~x[14] & x[55];
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & ~x[36] & ~x[42];
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & ~x[14];
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & x[55] & x[56];
			partial_clause[4][90] 	= partial_clause_prev[4][90] & ~x[14] & x[53] & x[54];
			partial_clause[4][91] 	= partial_clause_prev[4][91] & ~x[63];
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & ~x[18];
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & ~x[11];
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & ~x[13] & x[54] & x[55];
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & ~x[11];
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & ~x[0] & ~x[44];
			partial_clause[5][15] 	= partial_clause_prev[5][15] & x[60];
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & x[60];
			partial_clause[5][23] 	= partial_clause_prev[5][23] & ~x[41];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & ~x[44];
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & ~x[45];
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & ~x[45];
			partial_clause[5][50] 	= partial_clause_prev[5][50] & ~x[35] & ~x[62];
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & ~x[36] & ~x[63];
			partial_clause[5][55] 	= partial_clause_prev[5][55] & ~x[34] & ~x[62];
			partial_clause[5][56] 	= partial_clause_prev[5][56] & ~x[32];
			partial_clause[5][57] 	= partial_clause_prev[5][57] & ~x[63];
			partial_clause[5][58] 	= partial_clause_prev[5][58] & ~x[63];
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & ~x[34] & ~x[35] & ~x[39] & ~x[61];
			partial_clause[5][61] 	= partial_clause_prev[5][61] & ~x[15];
			partial_clause[5][62] 	= partial_clause_prev[5][62] & ~x[6];
			partial_clause[5][63] 	= partial_clause_prev[5][63] & ~x[61];
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & ~x[38] & ~x[63];
			partial_clause[5][66] 	= partial_clause_prev[5][66] & ~x[6] & ~x[35];
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & ~x[9] & ~x[34] & ~x[63];
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & ~x[39];
			partial_clause[5][72] 	= partial_clause_prev[5][72] & ~x[9] & ~x[34] & ~x[63];
			partial_clause[5][73] 	= partial_clause_prev[5][73] & ~x[7] & ~x[35] & ~x[61];
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & ~x[6] & ~x[33] & ~x[35] & ~x[63];
			partial_clause[5][76] 	= partial_clause_prev[5][76] & ~x[14] & ~x[63];
			partial_clause[5][77] 	= partial_clause_prev[5][77] & ~x[63];
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & ~x[36];
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & ~x[34];
			partial_clause[5][83] 	= partial_clause_prev[5][83] & ~x[34] & ~x[62];
			partial_clause[5][84] 	= partial_clause_prev[5][84] & ~x[63];
			partial_clause[5][85] 	= partial_clause_prev[5][85] & ~x[63];
			partial_clause[5][86] 	= partial_clause_prev[5][86] & ~x[8];
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & ~x[33];
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & ~x[63];
			partial_clause[5][93] 	= partial_clause_prev[5][93] & ~x[33] & ~x[34];
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & ~x[34];
			partial_clause[5][97] 	= partial_clause_prev[5][97] & ~x[63];
			partial_clause[5][98] 	= partial_clause_prev[5][98] & ~x[63];
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & ~x[37] & ~x[59];
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & ~x[11];
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & ~x[60];
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & ~x[62];
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & ~x[59];
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & ~x[61];
			partial_clause[6][34] 	= partial_clause_prev[6][34] & ~x[62];
			partial_clause[6][35] 	= partial_clause_prev[6][35] & ~x[46] & ~x[63];
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & ~x[61];
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & ~x[35];
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & ~x[3];
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & ~x[39];
			partial_clause[6][56] 	= partial_clause_prev[6][56] & ~x[7];
			partial_clause[6][57] 	= partial_clause_prev[6][57] & ~x[2] & ~x[4];
			partial_clause[6][58] 	= partial_clause_prev[6][58] & ~x[6];
			partial_clause[6][59] 	= partial_clause_prev[6][59] & ~x[41];
			partial_clause[6][60] 	= partial_clause_prev[6][60] & ~x[5];
			partial_clause[6][61] 	= partial_clause_prev[6][61] & ~x[3] & ~x[4] & ~x[6];
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & ~x[6];
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & ~x[3];
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & ~x[5];
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & ~x[35];
			partial_clause[6][72] 	= partial_clause_prev[6][72] & ~x[3];
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & ~x[5] & ~x[44];
			partial_clause[6][78] 	= partial_clause_prev[6][78] & ~x[5] & ~x[41];
			partial_clause[6][79] 	= partial_clause_prev[6][79] & ~x[2] & ~x[3];
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & ~x[5];
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & ~x[43];
			partial_clause[6][84] 	= partial_clause_prev[6][84] & ~x[3];
			partial_clause[6][85] 	= partial_clause_prev[6][85] & ~x[2] & ~x[3] & ~x[4];
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & ~x[5];
			partial_clause[6][89] 	= partial_clause_prev[6][89] & ~x[1] & ~x[4] & ~x[8];
			partial_clause[6][90] 	= partial_clause_prev[6][90] & ~x[7];
			partial_clause[6][91] 	= partial_clause_prev[6][91] & ~x[3];
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & ~x[4];
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & ~x[10];
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & ~x[5];
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & ~x[24] & ~x[26];
			partial_clause[7][2] 	= partial_clause_prev[7][2] & ~x[25] & ~x[26] & ~x[27] & ~x[29];
			partial_clause[7][3] 	= partial_clause_prev[7][3] & ~x[25] & ~x[28] & ~x[29];
			partial_clause[7][4] 	= partial_clause_prev[7][4] & ~x[9] & ~x[28];
			partial_clause[7][5] 	= partial_clause_prev[7][5] & ~x[22] & ~x[28] & ~x[31];
			partial_clause[7][6] 	= partial_clause_prev[7][6] & ~x[25] & ~x[28];
			partial_clause[7][7] 	= partial_clause_prev[7][7] & ~x[27] & ~x[28] & ~x[31];
			partial_clause[7][8] 	= partial_clause_prev[7][8] & ~x[23] & ~x[29];
			partial_clause[7][9] 	= partial_clause_prev[7][9] & ~x[25] & ~x[27] & ~x[33];
			partial_clause[7][10] 	= partial_clause_prev[7][10] & ~x[2] & ~x[25] & ~x[28];
			partial_clause[7][11] 	= partial_clause_prev[7][11] & ~x[23] & ~x[28];
			partial_clause[7][12] 	= partial_clause_prev[7][12] & ~x[25];
			partial_clause[7][13] 	= partial_clause_prev[7][13] & ~x[24] & ~x[28];
			partial_clause[7][14] 	= partial_clause_prev[7][14] & ~x[29] & ~x[32];
			partial_clause[7][15] 	= partial_clause_prev[7][15] & ~x[26] & ~x[27];
			partial_clause[7][16] 	= partial_clause_prev[7][16] & ~x[63];
			partial_clause[7][17] 	= partial_clause_prev[7][17] & ~x[0] & ~x[27] & ~x[30];
			partial_clause[7][18] 	= partial_clause_prev[7][18] & ~x[27];
			partial_clause[7][19] 	= partial_clause_prev[7][19] & ~x[25] & ~x[28] & ~x[29];
			partial_clause[7][20] 	= partial_clause_prev[7][20] & ~x[24] & ~x[27] & ~x[35];
			partial_clause[7][21] 	= partial_clause_prev[7][21] & ~x[26] & ~x[29] & ~x[30];
			partial_clause[7][22] 	= partial_clause_prev[7][22] & ~x[24] & ~x[28] & ~x[30];
			partial_clause[7][23] 	= partial_clause_prev[7][23] & ~x[13] & ~x[26] & ~x[28] & ~x[31];
			partial_clause[7][24] 	= partial_clause_prev[7][24] & ~x[4] & ~x[25] & ~x[26];
			partial_clause[7][25] 	= partial_clause_prev[7][25] & ~x[3];
			partial_clause[7][26] 	= partial_clause_prev[7][26] & ~x[29];
			partial_clause[7][27] 	= partial_clause_prev[7][27] & ~x[24] & ~x[29] & ~x[32];
			partial_clause[7][28] 	= partial_clause_prev[7][28] & ~x[0];
			partial_clause[7][29] 	= partial_clause_prev[7][29] & ~x[23] & ~x[26] & ~x[28];
			partial_clause[7][30] 	= partial_clause_prev[7][30] & ~x[25] & ~x[26];
			partial_clause[7][31] 	= partial_clause_prev[7][31] & ~x[28];
			partial_clause[7][32] 	= partial_clause_prev[7][32] & ~x[25] & ~x[27] & ~x[29] & ~x[62];
			partial_clause[7][33] 	= partial_clause_prev[7][33] & ~x[26] & ~x[28];
			partial_clause[7][34] 	= partial_clause_prev[7][34] & ~x[26] & ~x[62];
			partial_clause[7][35] 	= partial_clause_prev[7][35] & ~x[20] & ~x[21] & ~x[25] & ~x[31];
			partial_clause[7][36] 	= partial_clause_prev[7][36] & ~x[28] & ~x[32];
			partial_clause[7][37] 	= partial_clause_prev[7][37] & ~x[24] & ~x[26];
			partial_clause[7][38] 	= partial_clause_prev[7][38] & ~x[24] & ~x[28];
			partial_clause[7][39] 	= partial_clause_prev[7][39] & ~x[28];
			partial_clause[7][40] 	= partial_clause_prev[7][40] & ~x[24] & ~x[27];
			partial_clause[7][41] 	= partial_clause_prev[7][41] & ~x[29];
			partial_clause[7][42] 	= partial_clause_prev[7][42] & ~x[26];
			partial_clause[7][43] 	= partial_clause_prev[7][43] & ~x[3];
			partial_clause[7][44] 	= partial_clause_prev[7][44] & ~x[24] & ~x[27] & ~x[34];
			partial_clause[7][45] 	= partial_clause_prev[7][45] & ~x[27];
			partial_clause[7][46] 	= partial_clause_prev[7][46] & ~x[26] & ~x[27];
			partial_clause[7][47] 	= partial_clause_prev[7][47] & ~x[7] & ~x[27] & ~x[38];
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & ~x[2] & ~x[26];
			partial_clause[7][50] 	= partial_clause_prev[7][50] & x[27];
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & x[26] & ~x[42];
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & x[28];
			partial_clause[7][62] 	= partial_clause_prev[7][62] & x[57];
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & ~x[43];
			partial_clause[7][80] 	= partial_clause_prev[7][80] & x[55];
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & ~x[44];
			partial_clause[7][83] 	= partial_clause_prev[7][83] & x[28];
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & ~x[16];
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & ~x[14] & ~x[44];
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & ~x[44];
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & ~x[7];
			partial_clause[8][2] 	= partial_clause_prev[8][2] & ~x[16];
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & ~x[46];
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & ~x[16] & ~x[18];
			partial_clause[8][9] 	= partial_clause_prev[8][9] & ~x[46];
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & ~x[7];
			partial_clause[8][17] 	= partial_clause_prev[8][17] & ~x[20] & ~x[41];
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & ~x[45];
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & x[55];
			partial_clause[8][27] 	= partial_clause_prev[8][27] & ~x[7];
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & ~x[16];
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & ~x[12] & ~x[15] & ~x[19];
			partial_clause[8][33] 	= partial_clause_prev[8][33] & ~x[8];
			partial_clause[8][34] 	= partial_clause_prev[8][34] & x[28];
			partial_clause[8][35] 	= partial_clause_prev[8][35] & ~x[18] & ~x[45];
			partial_clause[8][36] 	= partial_clause_prev[8][36] & ~x[7];
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & ~x[19];
			partial_clause[8][40] 	= partial_clause_prev[8][40] & ~x[18];
			partial_clause[8][41] 	= partial_clause_prev[8][41] & ~x[17];
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & ~x[13];
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & ~x[41];
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & ~x[10];
			partial_clause[8][68] 	= partial_clause_prev[8][68] & ~x[42];
			partial_clause[8][69] 	= partial_clause_prev[8][69] & ~x[11];
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & ~x[44];
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & ~x[7];
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & ~x[14] & ~x[38];
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & ~x[26] & ~x[54];
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & ~x[9] & ~x[42];
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & ~x[16];
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & ~x[7];
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & ~x[43];
			partial_clause[8][94] 	= partial_clause_prev[8][94] & ~x[15];
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & ~x[53];
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & ~x[18] & ~x[30] & ~x[31];
			partial_clause[9][1] 	= partial_clause_prev[9][1] & ~x[28];
			partial_clause[9][2] 	= partial_clause_prev[9][2] & ~x[49];
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & ~x[26] & ~x[28];
			partial_clause[9][5] 	= partial_clause_prev[9][5] & ~x[25] & ~x[28] & ~x[31] & ~x[48] & ~x[62];
			partial_clause[9][6] 	= partial_clause_prev[9][6] & ~x[23] & ~x[28];
			partial_clause[9][7] 	= partial_clause_prev[9][7] & ~x[29];
			partial_clause[9][8] 	= partial_clause_prev[9][8] & ~x[49] & ~x[62];
			partial_clause[9][9] 	= partial_clause_prev[9][9] & ~x[13] & ~x[24] & ~x[27] & ~x[30];
			partial_clause[9][10] 	= partial_clause_prev[9][10] & ~x[26];
			partial_clause[9][11] 	= partial_clause_prev[9][11] & ~x[22] & ~x[27];
			partial_clause[9][12] 	= partial_clause_prev[9][12] & ~x[1] & ~x[3] & ~x[25];
			partial_clause[9][13] 	= partial_clause_prev[9][13] & ~x[31] & ~x[50];
			partial_clause[9][14] 	= partial_clause_prev[9][14] & ~x[25] & ~x[28] & ~x[30];
			partial_clause[9][15] 	= partial_clause_prev[9][15] & ~x[25] & ~x[27] & ~x[29] & ~x[32];
			partial_clause[9][16] 	= partial_clause_prev[9][16] & ~x[19] & ~x[24] & ~x[30];
			partial_clause[9][17] 	= partial_clause_prev[9][17] & ~x[31] & ~x[47] & ~x[48];
			partial_clause[9][18] 	= partial_clause_prev[9][18] & ~x[28];
			partial_clause[9][19] 	= partial_clause_prev[9][19] & ~x[25] & ~x[29];
			partial_clause[9][20] 	= partial_clause_prev[9][20] & ~x[1] & ~x[26];
			partial_clause[9][21] 	= partial_clause_prev[9][21] & ~x[50];
			partial_clause[9][22] 	= partial_clause_prev[9][22] & ~x[27];
			partial_clause[9][23] 	= partial_clause_prev[9][23] & ~x[22] & ~x[27] & ~x[29] & ~x[33] & ~x[62];
			partial_clause[9][24] 	= partial_clause_prev[9][24] & ~x[24] & ~x[26] & ~x[28] & ~x[48] & ~x[49];
			partial_clause[9][25] 	= partial_clause_prev[9][25] & ~x[1] & ~x[30];
			partial_clause[9][26] 	= partial_clause_prev[9][26] & ~x[26] & ~x[28] & ~x[29] & ~x[38] & ~x[63];
			partial_clause[9][27] 	= partial_clause_prev[9][27] & ~x[25] & ~x[30];
			partial_clause[9][28] 	= partial_clause_prev[9][28] & ~x[24] & ~x[63];
			partial_clause[9][29] 	= partial_clause_prev[9][29] & ~x[26] & ~x[29] & ~x[50];
			partial_clause[9][30] 	= partial_clause_prev[9][30] & ~x[26] & ~x[27] & ~x[29] & ~x[31] & ~x[45];
			partial_clause[9][31] 	= partial_clause_prev[9][31] & ~x[25] & ~x[28] & ~x[29] & ~x[50];
			partial_clause[9][32] 	= partial_clause_prev[9][32] & ~x[24] & ~x[50];
			partial_clause[9][33] 	= partial_clause_prev[9][33] & ~x[24] & ~x[27];
			partial_clause[9][34] 	= partial_clause_prev[9][34] & ~x[26] & ~x[28] & ~x[49] & ~x[61];
			partial_clause[9][35] 	= partial_clause_prev[9][35] & ~x[23] & ~x[29];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & ~x[0] & ~x[27] & ~x[29] & ~x[31];
			partial_clause[9][37] 	= partial_clause_prev[9][37] & ~x[28];
			partial_clause[9][38] 	= partial_clause_prev[9][38] & ~x[23];
			partial_clause[9][39] 	= partial_clause_prev[9][39] & ~x[27] & ~x[29];
			partial_clause[9][40] 	= partial_clause_prev[9][40] & ~x[25] & ~x[27] & ~x[29] & ~x[63];
			partial_clause[9][41] 	= partial_clause_prev[9][41] & ~x[27] & ~x[28] & ~x[30] & ~x[48];
			partial_clause[9][42] 	= partial_clause_prev[9][42] & ~x[27] & ~x[28] & ~x[30] & ~x[50];
			partial_clause[9][43] 	= partial_clause_prev[9][43] & ~x[30] & ~x[38] & ~x[62];
			partial_clause[9][44] 	= partial_clause_prev[9][44] & ~x[23] & ~x[29] & ~x[49];
			partial_clause[9][45] 	= partial_clause_prev[9][45] & ~x[18] & ~x[27] & ~x[28] & ~x[48];
			partial_clause[9][46] 	= partial_clause_prev[9][46] & ~x[26] & ~x[28] & ~x[29] & ~x[63];
			partial_clause[9][47] 	= partial_clause_prev[9][47] & ~x[24] & ~x[29] & ~x[31] & ~x[32];
			partial_clause[9][48] 	= partial_clause_prev[9][48] & ~x[28] & ~x[33] & ~x[36] & ~x[48] & ~x[61];
			partial_clause[9][49] 	= partial_clause_prev[9][49] & ~x[27] & ~x[49];
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & x[28];
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & x[28];
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & ~x[44];
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & ~x[16] & x[27];
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & x[29];
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & ~x[16];
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & x[25];
			partial_clause[9][91] 	= partial_clause_prev[9][91] & ~x[8];
			partial_clause[9][92] 	= partial_clause_prev[9][92] & ~x[7] & x[27] & ~x[42];
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & ~x[38];
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
		end
	end
endmodule


module HCB_3 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & ~x[10] & ~x[36] & ~x[63];
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & ~x[36] & ~x[58];
			partial_clause[0][8] 	= partial_clause_prev[0][8] & ~x[37];
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & ~x[7];
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & ~x[37] & ~x[63];
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & ~x[62];
			partial_clause[0][32] 	= partial_clause_prev[0][32] & ~x[57];
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & ~x[29];
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & ~x[62];
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & ~x[9];
			partial_clause[0][48] 	= partial_clause_prev[0][48] & ~x[58];
			partial_clause[0][49] 	= partial_clause_prev[0][49] & ~x[0];
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & ~x[4];
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & ~x[32];
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & ~x[56];
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & ~x[31];
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & ~x[3];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & ~x[4] & ~x[59];
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & ~x[60];
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & ~x[58];
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & ~x[59];
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & ~x[3] & ~x[7] & ~x[62];
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & ~x[2];
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & ~x[2];
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & ~x[62];
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & ~x[39];
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & ~x[14];
			partial_clause[1][4] 	= partial_clause_prev[1][4] & ~x[42];
			partial_clause[1][5] 	= partial_clause_prev[1][5] & ~x[41];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & ~x[40];
			partial_clause[1][7] 	= partial_clause_prev[1][7] & ~x[26] & ~x[33];
			partial_clause[1][8] 	= partial_clause_prev[1][8] & ~x[14];
			partial_clause[1][9] 	= partial_clause_prev[1][9] & ~x[13];
			partial_clause[1][10] 	= partial_clause_prev[1][10] & ~x[43];
			partial_clause[1][11] 	= partial_clause_prev[1][11] & ~x[40];
			partial_clause[1][12] 	= partial_clause_prev[1][12] & ~x[14] & ~x[40];
			partial_clause[1][13] 	= partial_clause_prev[1][13] & ~x[42];
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & ~x[14] & ~x[62];
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & ~x[14] & ~x[43];
			partial_clause[1][19] 	= partial_clause_prev[1][19] & ~x[42];
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & ~x[14];
			partial_clause[1][22] 	= partial_clause_prev[1][22] & ~x[42];
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & ~x[42];
			partial_clause[1][25] 	= partial_clause_prev[1][25] & ~x[14];
			partial_clause[1][26] 	= partial_clause_prev[1][26] & ~x[14];
			partial_clause[1][27] 	= partial_clause_prev[1][27] & ~x[14];
			partial_clause[1][28] 	= partial_clause_prev[1][28] & ~x[13] & ~x[42];
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & ~x[14];
			partial_clause[1][31] 	= partial_clause_prev[1][31] & ~x[42];
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & ~x[14] & ~x[41];
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & ~x[13];
			partial_clause[1][36] 	= partial_clause_prev[1][36] & ~x[13];
			partial_clause[1][37] 	= partial_clause_prev[1][37] & ~x[14] & ~x[54];
			partial_clause[1][38] 	= partial_clause_prev[1][38] & ~x[14];
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & ~x[15] & ~x[43];
			partial_clause[1][41] 	= partial_clause_prev[1][41] & ~x[52];
			partial_clause[1][42] 	= partial_clause_prev[1][42] & ~x[42];
			partial_clause[1][43] 	= partial_clause_prev[1][43] & ~x[43];
			partial_clause[1][44] 	= partial_clause_prev[1][44] & ~x[42];
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & ~x[41];
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & ~x[61];
			partial_clause[1][58] 	= partial_clause_prev[1][58] & ~x[60];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & ~x[59];
			partial_clause[1][65] 	= partial_clause_prev[1][65] & ~x[3];
			partial_clause[1][66] 	= partial_clause_prev[1][66] & ~x[34] & ~x[58];
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & ~x[2];
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & ~x[33];
			partial_clause[1][72] 	= partial_clause_prev[1][72] & ~x[32];
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & 1'b1;
			partial_clause[1][75] 	= partial_clause_prev[1][75] & ~x[6] & ~x[32];
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & ~x[63];
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & ~x[31];
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & ~x[62];
			partial_clause[1][82] 	= partial_clause_prev[1][82] & x[42];
			partial_clause[1][83] 	= partial_clause_prev[1][83] & ~x[34];
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & ~x[60] & ~x[61];
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & ~x[6];
			partial_clause[1][92] 	= partial_clause_prev[1][92] & ~x[6] & x[52] & ~x[61];
			partial_clause[1][93] 	= partial_clause_prev[1][93] & ~x[6];
			partial_clause[1][94] 	= partial_clause_prev[1][94] & ~x[4] & ~x[30] & ~x[32];
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & ~x[61];
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & ~x[63];
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & ~x[0];
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & ~x[35];
			partial_clause[2][13] 	= partial_clause_prev[2][13] & ~x[57];
			partial_clause[2][14] 	= partial_clause_prev[2][14] & ~x[7];
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & ~x[56];
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & ~x[29];
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & ~x[60];
			partial_clause[2][35] 	= partial_clause_prev[2][35] & ~x[30];
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & ~x[58];
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & ~x[27];
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & ~x[31];
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & ~x[10];
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & ~x[7];
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & 1'b1;
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & ~x[7];
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & ~x[9];
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & ~x[59];
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & ~x[58];
			partial_clause[2][92] 	= partial_clause_prev[2][92] & ~x[2];
			partial_clause[2][93] 	= partial_clause_prev[2][93] & ~x[4];
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & ~x[27] & ~x[56];
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & ~x[27];
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & ~x[28];
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & ~x[32];
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & ~x[55];
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & ~x[29];
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & ~x[27];
			partial_clause[3][29] 	= partial_clause_prev[3][29] & ~x[27];
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & ~x[56];
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & ~x[59];
			partial_clause[3][37] 	= partial_clause_prev[3][37] & ~x[56];
			partial_clause[3][38] 	= partial_clause_prev[3][38] & ~x[0] & ~x[27];
			partial_clause[3][39] 	= partial_clause_prev[3][39] & ~x[28];
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & ~x[1];
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & ~x[62];
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & ~x[10];
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & ~x[4];
			partial_clause[3][58] 	= partial_clause_prev[3][58] & ~x[32];
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & ~x[11];
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & ~x[9];
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[12];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & ~x[6];
			partial_clause[3][70] 	= partial_clause_prev[3][70] & ~x[11];
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & ~x[4];
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & ~x[2];
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & ~x[32];
			partial_clause[3][79] 	= partial_clause_prev[3][79] & ~x[13];
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & ~x[9];
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & ~x[35];
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & ~x[10];
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & ~x[8] & ~x[58];
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & ~x[8] & ~x[14];
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & ~x[20] & ~x[48];
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & ~x[19];
			partial_clause[4][4] 	= partial_clause_prev[4][4] & ~x[46];
			partial_clause[4][5] 	= partial_clause_prev[4][5] & ~x[47];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & ~x[19];
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & ~x[1] & ~x[47];
			partial_clause[4][9] 	= partial_clause_prev[4][9] & ~x[18];
			partial_clause[4][10] 	= partial_clause_prev[4][10] & ~x[47];
			partial_clause[4][11] 	= partial_clause_prev[4][11] & ~x[19] & ~x[47];
			partial_clause[4][12] 	= partial_clause_prev[4][12] & ~x[18];
			partial_clause[4][13] 	= partial_clause_prev[4][13] & ~x[18] & ~x[46];
			partial_clause[4][14] 	= partial_clause_prev[4][14] & ~x[18];
			partial_clause[4][15] 	= partial_clause_prev[4][15] & ~x[46];
			partial_clause[4][16] 	= partial_clause_prev[4][16] & ~x[47];
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & ~x[18] & ~x[46];
			partial_clause[4][20] 	= partial_clause_prev[4][20] & ~x[19] & ~x[47];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & ~x[47];
			partial_clause[4][22] 	= partial_clause_prev[4][22] & ~x[19];
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & ~x[19];
			partial_clause[4][25] 	= partial_clause_prev[4][25] & ~x[47];
			partial_clause[4][26] 	= partial_clause_prev[4][26] & ~x[46];
			partial_clause[4][27] 	= partial_clause_prev[4][27] & ~x[18] & ~x[46];
			partial_clause[4][28] 	= partial_clause_prev[4][28] & ~x[19];
			partial_clause[4][29] 	= partial_clause_prev[4][29] & ~x[47];
			partial_clause[4][30] 	= partial_clause_prev[4][30] & ~x[4] & ~x[19];
			partial_clause[4][31] 	= partial_clause_prev[4][31] & ~x[47];
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[5] & ~x[18];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & ~x[19];
			partial_clause[4][34] 	= partial_clause_prev[4][34] & ~x[17];
			partial_clause[4][35] 	= partial_clause_prev[4][35] & ~x[47];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & ~x[19];
			partial_clause[4][37] 	= partial_clause_prev[4][37] & ~x[18];
			partial_clause[4][38] 	= partial_clause_prev[4][38] & ~x[19] & ~x[47];
			partial_clause[4][39] 	= partial_clause_prev[4][39] & ~x[18];
			partial_clause[4][40] 	= partial_clause_prev[4][40] & ~x[47];
			partial_clause[4][41] 	= partial_clause_prev[4][41] & ~x[47];
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & ~x[19];
			partial_clause[4][46] 	= partial_clause_prev[4][46] & ~x[20] & ~x[48];
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & ~x[18];
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[19];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & x[20];
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & ~x[6];
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & x[19];
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & ~x[62];
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & x[16] & x[19];
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & x[19];
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & x[20] & ~x[31];
			partial_clause[4][74] 	= partial_clause_prev[4][74] & x[17] & ~x[60];
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & ~x[61];
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & ~x[59];
			partial_clause[4][86] 	= partial_clause_prev[4][86] & ~x[1] & x[45] & x[47] & ~x[61];
			partial_clause[4][87] 	= partial_clause_prev[4][87] & x[18] & x[19] & x[20];
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & ~x[62];
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & ~x[33];
			partial_clause[4][96] 	= partial_clause_prev[4][96] & ~x[29];
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & ~x[61];
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & x[56];
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & ~x[7];
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & x[56];
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & x[24];
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & ~x[55];
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & ~x[56] & ~x[60];
			partial_clause[5][53] 	= partial_clause_prev[5][53] & ~x[0] & ~x[28] & ~x[56];
			partial_clause[5][54] 	= partial_clause_prev[5][54] & ~x[29] & ~x[56];
			partial_clause[5][55] 	= partial_clause_prev[5][55] & ~x[28] & ~x[55];
			partial_clause[5][56] 	= partial_clause_prev[5][56] & ~x[56];
			partial_clause[5][57] 	= partial_clause_prev[5][57] & ~x[55];
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & ~x[31];
			partial_clause[5][60] 	= partial_clause_prev[5][60] & ~x[56];
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & ~x[4] & ~x[27] & ~x[57];
			partial_clause[5][63] 	= partial_clause_prev[5][63] & ~x[26] & ~x[58];
			partial_clause[5][64] 	= partial_clause_prev[5][64] & ~x[27];
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & ~x[27] & ~x[56];
			partial_clause[5][67] 	= partial_clause_prev[5][67] & ~x[0] & ~x[27] & ~x[28] & ~x[55];
			partial_clause[5][68] 	= partial_clause_prev[5][68] & ~x[55] & ~x[56];
			partial_clause[5][69] 	= partial_clause_prev[5][69] & ~x[29] & ~x[56];
			partial_clause[5][70] 	= partial_clause_prev[5][70] & ~x[26];
			partial_clause[5][71] 	= partial_clause_prev[5][71] & ~x[5] & ~x[28];
			partial_clause[5][72] 	= partial_clause_prev[5][72] & ~x[29] & ~x[34] & ~x[58];
			partial_clause[5][73] 	= partial_clause_prev[5][73] & ~x[26] & ~x[27];
			partial_clause[5][74] 	= partial_clause_prev[5][74] & ~x[28] & ~x[55] & ~x[56] & ~x[57];
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & ~x[27] & ~x[55];
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & ~x[2] & ~x[27] & ~x[57];
			partial_clause[5][79] 	= partial_clause_prev[5][79] & ~x[0] & ~x[27];
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & ~x[4] & ~x[27];
			partial_clause[5][83] 	= partial_clause_prev[5][83] & ~x[27] & ~x[28] & ~x[56];
			partial_clause[5][84] 	= partial_clause_prev[5][84] & ~x[55];
			partial_clause[5][85] 	= partial_clause_prev[5][85] & ~x[29] & ~x[55];
			partial_clause[5][86] 	= partial_clause_prev[5][86] & ~x[33];
			partial_clause[5][87] 	= partial_clause_prev[5][87] & ~x[28] & ~x[54];
			partial_clause[5][88] 	= partial_clause_prev[5][88] & ~x[26] & ~x[53];
			partial_clause[5][89] 	= partial_clause_prev[5][89] & ~x[55];
			partial_clause[5][90] 	= partial_clause_prev[5][90] & ~x[56] & ~x[57];
			partial_clause[5][91] 	= partial_clause_prev[5][91] & ~x[55];
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & ~x[0] & ~x[54];
			partial_clause[5][94] 	= partial_clause_prev[5][94] & ~x[0] & ~x[29];
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & ~x[27] & ~x[56];
			partial_clause[5][97] 	= partial_clause_prev[5][97] & ~x[59];
			partial_clause[5][98] 	= partial_clause_prev[5][98] & ~x[3] & ~x[27] & ~x[28] & ~x[57];
			partial_clause[5][99] 	= partial_clause_prev[5][99] & ~x[27];
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & ~x[23] & ~x[27] & ~x[52];
			partial_clause[6][1] 	= partial_clause_prev[6][1] & ~x[52];
			partial_clause[6][2] 	= partial_clause_prev[6][2] & ~x[51];
			partial_clause[6][3] 	= partial_clause_prev[6][3] & ~x[50];
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & ~x[51];
			partial_clause[6][6] 	= partial_clause_prev[6][6] & ~x[28] & ~x[51] & ~x[52];
			partial_clause[6][7] 	= partial_clause_prev[6][7] & ~x[53] & ~x[63];
			partial_clause[6][8] 	= partial_clause_prev[6][8] & ~x[50];
			partial_clause[6][9] 	= partial_clause_prev[6][9] & ~x[24];
			partial_clause[6][10] 	= partial_clause_prev[6][10] & ~x[23] & ~x[50] & ~x[52];
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & ~x[24];
			partial_clause[6][13] 	= partial_clause_prev[6][13] & ~x[23] & ~x[52];
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & ~x[26] & ~x[50];
			partial_clause[6][16] 	= partial_clause_prev[6][16] & ~x[24] & ~x[50];
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & ~x[52];
			partial_clause[6][19] 	= partial_clause_prev[6][19] & ~x[24];
			partial_clause[6][20] 	= partial_clause_prev[6][20] & ~x[51];
			partial_clause[6][21] 	= partial_clause_prev[6][21] & ~x[24] & ~x[51];
			partial_clause[6][22] 	= partial_clause_prev[6][22] & ~x[50] & ~x[51];
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & ~x[51];
			partial_clause[6][25] 	= partial_clause_prev[6][25] & ~x[10] & ~x[24] & ~x[54] & ~x[62];
			partial_clause[6][26] 	= partial_clause_prev[6][26] & ~x[52];
			partial_clause[6][27] 	= partial_clause_prev[6][27] & ~x[49] & ~x[51];
			partial_clause[6][28] 	= partial_clause_prev[6][28] & ~x[50] & ~x[52];
			partial_clause[6][29] 	= partial_clause_prev[6][29] & ~x[51];
			partial_clause[6][30] 	= partial_clause_prev[6][30] & ~x[23] & ~x[52] & ~x[53];
			partial_clause[6][31] 	= partial_clause_prev[6][31] & ~x[22] & ~x[48] & ~x[53];
			partial_clause[6][32] 	= partial_clause_prev[6][32] & ~x[51];
			partial_clause[6][33] 	= partial_clause_prev[6][33] & ~x[50];
			partial_clause[6][34] 	= partial_clause_prev[6][34] & ~x[23] & ~x[50] & ~x[51];
			partial_clause[6][35] 	= partial_clause_prev[6][35] & ~x[52];
			partial_clause[6][36] 	= partial_clause_prev[6][36] & ~x[52];
			partial_clause[6][37] 	= partial_clause_prev[6][37] & ~x[50] & ~x[51];
			partial_clause[6][38] 	= partial_clause_prev[6][38] & ~x[24] & ~x[51];
			partial_clause[6][39] 	= partial_clause_prev[6][39] & ~x[51] & ~x[53];
			partial_clause[6][40] 	= partial_clause_prev[6][40] & ~x[24] & ~x[37];
			partial_clause[6][41] 	= partial_clause_prev[6][41] & ~x[23] & ~x[50];
			partial_clause[6][42] 	= partial_clause_prev[6][42] & ~x[50] & ~x[56];
			partial_clause[6][43] 	= partial_clause_prev[6][43] & ~x[24];
			partial_clause[6][44] 	= partial_clause_prev[6][44] & ~x[24] & ~x[54];
			partial_clause[6][45] 	= partial_clause_prev[6][45] & ~x[2] & ~x[51];
			partial_clause[6][46] 	= partial_clause_prev[6][46] & ~x[23] & ~x[50] & ~x[51] & ~x[53];
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & ~x[27] & ~x[37];
			partial_clause[6][49] 	= partial_clause_prev[6][49] & ~x[30] & ~x[50] & ~x[52];
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & x[51];
			partial_clause[6][53] 	= partial_clause_prev[6][53] & x[51] & ~x[59];
			partial_clause[6][54] 	= partial_clause_prev[6][54] & ~x[61];
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & x[50];
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & ~x[30] & ~x[35];
			partial_clause[6][71] 	= partial_clause_prev[6][71] & x[22];
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & ~x[61];
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & x[51];
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & ~x[5] & x[23];
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & ~x[59];
			partial_clause[6][91] 	= partial_clause_prev[6][91] & ~x[31];
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & ~x[30];
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & ~x[31];
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & ~x[0];
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & ~x[0];
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & ~x[38];
			partial_clause[7][55] 	= partial_clause_prev[7][55] & ~x[38];
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & ~x[38];
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & ~x[7];
			partial_clause[7][60] 	= partial_clause_prev[7][60] & ~x[38];
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & ~x[9];
			partial_clause[7][63] 	= partial_clause_prev[7][63] & ~x[30];
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & ~x[62];
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & ~x[3] & ~x[61];
			partial_clause[7][83] 	= partial_clause_prev[7][83] & ~x[8] & ~x[37];
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & ~x[8];
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & ~x[39];
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & ~x[38];
			partial_clause[7][96] 	= partial_clause_prev[7][96] & ~x[38];
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & ~x[63];
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & ~x[63];
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & ~x[8];
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & ~x[2] & ~x[36];
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & ~x[8] & ~x[61];
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & ~x[8];
			partial_clause[8][17] 	= partial_clause_prev[8][17] & ~x[63];
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & ~x[8];
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & ~x[37];
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & ~x[7];
			partial_clause[8][44] 	= partial_clause_prev[8][44] & ~x[9];
			partial_clause[8][45] 	= partial_clause_prev[8][45] & ~x[5];
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & ~x[60];
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & ~x[3];
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & ~x[31] & ~x[56];
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & ~x[61];
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & ~x[3] & ~x[54];
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & ~x[56];
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & ~x[31];
			partial_clause[8][68] 	= partial_clause_prev[8][68] & ~x[4];
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & ~x[62];
			partial_clause[8][74] 	= partial_clause_prev[8][74] & ~x[1];
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & ~x[59];
			partial_clause[8][77] 	= partial_clause_prev[8][77] & ~x[3];
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & ~x[28] & ~x[56];
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & ~x[2] & ~x[55];
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & ~x[2] & ~x[28] & ~x[59];
			partial_clause[8][88] 	= partial_clause_prev[8][88] & ~x[28] & ~x[33];
			partial_clause[8][89] 	= partial_clause_prev[8][89] & ~x[56];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & ~x[26];
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & ~x[3] & ~x[26];
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & ~x[39] & ~x[55];
			partial_clause[9][1] 	= partial_clause_prev[9][1] & x[19] & ~x[39];
			partial_clause[9][2] 	= partial_clause_prev[9][2] & x[19] & ~x[39];
			partial_clause[9][3] 	= partial_clause_prev[9][3] & ~x[7] & ~x[10] & x[19] & ~x[26];
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & x[20];
			partial_clause[9][7] 	= partial_clause_prev[9][7] & ~x[12];
			partial_clause[9][8] 	= partial_clause_prev[9][8] & ~x[13] & x[19] & x[20];
			partial_clause[9][9] 	= partial_clause_prev[9][9] & x[18] & x[19] & ~x[27] & ~x[39];
			partial_clause[9][10] 	= partial_clause_prev[9][10] & x[18];
			partial_clause[9][11] 	= partial_clause_prev[9][11] & x[18] & ~x[26];
			partial_clause[9][12] 	= partial_clause_prev[9][12] & x[19] & ~x[39];
			partial_clause[9][13] 	= partial_clause_prev[9][13] & x[19];
			partial_clause[9][14] 	= partial_clause_prev[9][14] & x[19];
			partial_clause[9][15] 	= partial_clause_prev[9][15] & ~x[27];
			partial_clause[9][16] 	= partial_clause_prev[9][16] & ~x[11] & x[17];
			partial_clause[9][17] 	= partial_clause_prev[9][17] & x[19] & ~x[27] & ~x[37];
			partial_clause[9][18] 	= partial_clause_prev[9][18] & ~x[12] & x[19];
			partial_clause[9][19] 	= partial_clause_prev[9][19] & x[18];
			partial_clause[9][20] 	= partial_clause_prev[9][20] & x[19];
			partial_clause[9][21] 	= partial_clause_prev[9][21] & ~x[13] & x[19];
			partial_clause[9][22] 	= partial_clause_prev[9][22] & x[19];
			partial_clause[9][23] 	= partial_clause_prev[9][23] & ~x[12] & ~x[37];
			partial_clause[9][24] 	= partial_clause_prev[9][24] & x[19] & ~x[39];
			partial_clause[9][25] 	= partial_clause_prev[9][25] & ~x[12] & x[20];
			partial_clause[9][26] 	= partial_clause_prev[9][26] & x[19] & ~x[27];
			partial_clause[9][27] 	= partial_clause_prev[9][27] & x[18];
			partial_clause[9][28] 	= partial_clause_prev[9][28] & x[18] & ~x[26] & ~x[37];
			partial_clause[9][29] 	= partial_clause_prev[9][29] & x[19] & ~x[38] & ~x[63];
			partial_clause[9][30] 	= partial_clause_prev[9][30] & ~x[11] & x[18];
			partial_clause[9][31] 	= partial_clause_prev[9][31] & ~x[12] & ~x[26];
			partial_clause[9][32] 	= partial_clause_prev[9][32] & x[19] & ~x[39];
			partial_clause[9][33] 	= partial_clause_prev[9][33] & ~x[12] & x[18] & ~x[38];
			partial_clause[9][34] 	= partial_clause_prev[9][34] & x[18] & x[19];
			partial_clause[9][35] 	= partial_clause_prev[9][35] & ~x[12];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & ~x[12] & x[20];
			partial_clause[9][37] 	= partial_clause_prev[9][37] & x[20] & ~x[39];
			partial_clause[9][38] 	= partial_clause_prev[9][38] & ~x[9] & x[18] & ~x[26] & ~x[37];
			partial_clause[9][39] 	= partial_clause_prev[9][39] & x[20];
			partial_clause[9][40] 	= partial_clause_prev[9][40] & ~x[11] & x[19] & ~x[39] & ~x[55];
			partial_clause[9][41] 	= partial_clause_prev[9][41] & x[19];
			partial_clause[9][42] 	= partial_clause_prev[9][42] & x[19] & ~x[27];
			partial_clause[9][43] 	= partial_clause_prev[9][43] & x[19];
			partial_clause[9][44] 	= partial_clause_prev[9][44] & x[20] & ~x[39];
			partial_clause[9][45] 	= partial_clause_prev[9][45] & x[19];
			partial_clause[9][46] 	= partial_clause_prev[9][46] & ~x[12] & x[19] & x[46];
			partial_clause[9][47] 	= partial_clause_prev[9][47] & ~x[26];
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & ~x[12] & x[19] & ~x[27];
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & ~x[7];
			partial_clause[9][54] 	= partial_clause_prev[9][54] & ~x[58];
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & ~x[6];
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & ~x[1];
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & ~x[20];
			partial_clause[9][70] 	= partial_clause_prev[9][70] & ~x[30];
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & ~x[0] & ~x[28];
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
		end
	end
endmodule


module HCB_4 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & ~x[1] & ~x[54];
			partial_clause[0][3] 	= partial_clause_prev[0][3] & ~x[21];
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & ~x[55];
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & ~x[26] & ~x[51];
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & ~x[56];
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & ~x[27];
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & ~x[25] & ~x[26] & ~x[28];
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & ~x[0];
			partial_clause[0][41] 	= partial_clause_prev[0][41] & ~x[27] & ~x[51];
			partial_clause[0][42] 	= partial_clause_prev[0][42] & ~x[28];
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & ~x[55];
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & ~x[0] & ~x[25];
			partial_clause[0][50] 	= partial_clause_prev[0][50] & ~x[51];
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & ~x[24];
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & ~x[54];
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & ~x[53];
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & ~x[53];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & ~x[24];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & ~x[48];
			partial_clause[0][75] 	= partial_clause_prev[0][75] & ~x[24];
			partial_clause[0][76] 	= partial_clause_prev[0][76] & ~x[22] & ~x[53];
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & ~x[54];
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & ~x[50];
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & ~x[53];
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & ~x[23];
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & ~x[54];
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & ~x[56];
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[34] & ~x[46];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & ~x[63];
			partial_clause[1][2] 	= partial_clause_prev[1][2] & ~x[7] & ~x[22] & ~x[44] & ~x[63];
			partial_clause[1][3] 	= partial_clause_prev[1][3] & ~x[35];
			partial_clause[1][4] 	= partial_clause_prev[1][4] & ~x[63];
			partial_clause[1][5] 	= partial_clause_prev[1][5] & ~x[44];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & ~x[16];
			partial_clause[1][7] 	= partial_clause_prev[1][7] & ~x[2];
			partial_clause[1][8] 	= partial_clause_prev[1][8] & ~x[34] & ~x[46];
			partial_clause[1][9] 	= partial_clause_prev[1][9] & ~x[34];
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & ~x[34] & ~x[62];
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & ~x[6] & ~x[34];
			partial_clause[1][15] 	= partial_clause_prev[1][15] & ~x[15] & ~x[35];
			partial_clause[1][16] 	= partial_clause_prev[1][16] & ~x[7] & ~x[63];
			partial_clause[1][17] 	= partial_clause_prev[1][17] & ~x[7];
			partial_clause[1][18] 	= partial_clause_prev[1][18] & ~x[18] & ~x[34];
			partial_clause[1][19] 	= partial_clause_prev[1][19] & ~x[20] & ~x[35];
			partial_clause[1][20] 	= partial_clause_prev[1][20] & ~x[4];
			partial_clause[1][21] 	= partial_clause_prev[1][21] & ~x[7];
			partial_clause[1][22] 	= partial_clause_prev[1][22] & ~x[7] & x[39] & ~x[45];
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & ~x[63];
			partial_clause[1][25] 	= partial_clause_prev[1][25] & ~x[6] & ~x[45];
			partial_clause[1][26] 	= partial_clause_prev[1][26] & ~x[45] & ~x[63];
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & ~x[63];
			partial_clause[1][29] 	= partial_clause_prev[1][29] & ~x[5] & ~x[17] & ~x[61];
			partial_clause[1][30] 	= partial_clause_prev[1][30] & ~x[17];
			partial_clause[1][31] 	= partial_clause_prev[1][31] & ~x[63];
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & ~x[43] & ~x[63];
			partial_clause[1][34] 	= partial_clause_prev[1][34] & ~x[7] & ~x[35] & ~x[63];
			partial_clause[1][35] 	= partial_clause_prev[1][35] & ~x[17] & ~x[63];
			partial_clause[1][36] 	= partial_clause_prev[1][36] & ~x[1] & ~x[6];
			partial_clause[1][37] 	= partial_clause_prev[1][37] & ~x[63];
			partial_clause[1][38] 	= partial_clause_prev[1][38] & ~x[34];
			partial_clause[1][39] 	= partial_clause_prev[1][39] & ~x[60];
			partial_clause[1][40] 	= partial_clause_prev[1][40] & ~x[57];
			partial_clause[1][41] 	= partial_clause_prev[1][41] & ~x[6];
			partial_clause[1][42] 	= partial_clause_prev[1][42] & ~x[35];
			partial_clause[1][43] 	= partial_clause_prev[1][43] & ~x[18] & ~x[63];
			partial_clause[1][44] 	= partial_clause_prev[1][44] & ~x[5] & ~x[6];
			partial_clause[1][45] 	= partial_clause_prev[1][45] & ~x[63];
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & ~x[6] & ~x[18];
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & ~x[5] & ~x[32];
			partial_clause[1][50] 	= partial_clause_prev[1][50] & ~x[50];
			partial_clause[1][51] 	= partial_clause_prev[1][51] & ~x[22];
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & x[7] & ~x[52];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & x[7];
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & x[61];
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & ~x[24];
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & ~x[53] & ~x[54];
			partial_clause[1][69] 	= partial_clause_prev[1][69] & ~x[53];
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & x[7];
			partial_clause[1][72] 	= partial_clause_prev[1][72] & x[61];
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & 1'b1;
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & ~x[23];
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & ~x[52];
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & x[6] & ~x[26];
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & ~x[22];
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & ~x[50] & ~x[54];
			partial_clause[1][91] 	= partial_clause_prev[1][91] & ~x[24];
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & x[62];
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & ~x[54] & x[63];
			partial_clause[1][98] 	= partial_clause_prev[1][98] & x[6] & ~x[23];
			partial_clause[1][99] 	= partial_clause_prev[1][99] & ~x[53];
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & ~x[55];
			partial_clause[2][1] 	= partial_clause_prev[2][1] & ~x[28];
			partial_clause[2][2] 	= partial_clause_prev[2][2] & ~x[27];
			partial_clause[2][3] 	= partial_clause_prev[2][3] & ~x[60] & ~x[63];
			partial_clause[2][4] 	= partial_clause_prev[2][4] & ~x[63];
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & ~x[48] & ~x[54];
			partial_clause[2][7] 	= partial_clause_prev[2][7] & ~x[60];
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & ~x[20] & ~x[61] & ~x[63];
			partial_clause[2][11] 	= partial_clause_prev[2][11] & ~x[20];
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & ~x[63];
			partial_clause[2][17] 	= partial_clause_prev[2][17] & ~x[61] & ~x[63];
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & ~x[61];
			partial_clause[2][28] 	= partial_clause_prev[2][28] & ~x[63];
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & ~x[63];
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & ~x[59];
			partial_clause[2][34] 	= partial_clause_prev[2][34] & ~x[60];
			partial_clause[2][35] 	= partial_clause_prev[2][35] & ~x[62];
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & ~x[61];
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & ~x[38];
			partial_clause[2][40] 	= partial_clause_prev[2][40] & ~x[63];
			partial_clause[2][41] 	= partial_clause_prev[2][41] & ~x[37];
			partial_clause[2][42] 	= partial_clause_prev[2][42] & ~x[60] & ~x[62];
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & ~x[60];
			partial_clause[2][45] 	= partial_clause_prev[2][45] & ~x[53] & ~x[62];
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & ~x[49];
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & ~x[52];
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & ~x[51];
			partial_clause[2][56] 	= partial_clause_prev[2][56] & ~x[51];
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & x[63];
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & ~x[23];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & ~x[50];
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & ~x[50];
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & ~x[53];
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & x[63];
			partial_clause[2][99] 	= partial_clause_prev[2][99] & ~x[23] & ~x[27];
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & ~x[7];
			partial_clause[3][1] 	= partial_clause_prev[3][1] & ~x[22];
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & ~x[32] & ~x[57];
			partial_clause[3][5] 	= partial_clause_prev[3][5] & ~x[34] & ~x[35] & ~x[60];
			partial_clause[3][6] 	= partial_clause_prev[3][6] & ~x[23] & ~x[59] & ~x[60];
			partial_clause[3][7] 	= partial_clause_prev[3][7] & ~x[60];
			partial_clause[3][8] 	= partial_clause_prev[3][8] & ~x[26] & ~x[35] & ~x[61];
			partial_clause[3][9] 	= partial_clause_prev[3][9] & ~x[33] & ~x[34] & ~x[59];
			partial_clause[3][10] 	= partial_clause_prev[3][10] & ~x[34] & ~x[57];
			partial_clause[3][11] 	= partial_clause_prev[3][11] & ~x[20] & ~x[34];
			partial_clause[3][12] 	= partial_clause_prev[3][12] & ~x[60] & ~x[62];
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & ~x[19] & ~x[34] & ~x[58];
			partial_clause[3][15] 	= partial_clause_prev[3][15] & ~x[34];
			partial_clause[3][16] 	= partial_clause_prev[3][16] & ~x[62];
			partial_clause[3][17] 	= partial_clause_prev[3][17] & ~x[35] & ~x[61];
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & ~x[35] & ~x[60];
			partial_clause[3][20] 	= partial_clause_prev[3][20] & ~x[34] & ~x[59];
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & ~x[35] & ~x[59];
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & ~x[35] & ~x[61];
			partial_clause[3][25] 	= partial_clause_prev[3][25] & ~x[58] & ~x[60];
			partial_clause[3][26] 	= partial_clause_prev[3][26] & ~x[48] & ~x[51] & ~x[60] & ~x[61];
			partial_clause[3][27] 	= partial_clause_prev[3][27] & ~x[34] & ~x[47];
			partial_clause[3][28] 	= partial_clause_prev[3][28] & ~x[34];
			partial_clause[3][29] 	= partial_clause_prev[3][29] & ~x[8] & ~x[59] & ~x[60];
			partial_clause[3][30] 	= partial_clause_prev[3][30] & ~x[35] & ~x[60];
			partial_clause[3][31] 	= partial_clause_prev[3][31] & ~x[33] & ~x[34];
			partial_clause[3][32] 	= partial_clause_prev[3][32] & ~x[34] & ~x[60];
			partial_clause[3][33] 	= partial_clause_prev[3][33] & ~x[33];
			partial_clause[3][34] 	= partial_clause_prev[3][34] & ~x[34];
			partial_clause[3][35] 	= partial_clause_prev[3][35] & ~x[35] & ~x[61];
			partial_clause[3][36] 	= partial_clause_prev[3][36] & ~x[60];
			partial_clause[3][37] 	= partial_clause_prev[3][37] & ~x[34] & ~x[59] & ~x[60];
			partial_clause[3][38] 	= partial_clause_prev[3][38] & ~x[60];
			partial_clause[3][39] 	= partial_clause_prev[3][39] & ~x[34] & ~x[60];
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & ~x[22] & ~x[35] & ~x[60];
			partial_clause[3][42] 	= partial_clause_prev[3][42] & ~x[32];
			partial_clause[3][43] 	= partial_clause_prev[3][43] & ~x[60] & ~x[61];
			partial_clause[3][44] 	= partial_clause_prev[3][44] & ~x[21] & ~x[34] & ~x[35] & ~x[46] & ~x[61];
			partial_clause[3][45] 	= partial_clause_prev[3][45] & ~x[32] & ~x[50];
			partial_clause[3][46] 	= partial_clause_prev[3][46] & ~x[25] & ~x[35];
			partial_clause[3][47] 	= partial_clause_prev[3][47] & ~x[53];
			partial_clause[3][48] 	= partial_clause_prev[3][48] & ~x[35] & ~x[60];
			partial_clause[3][49] 	= partial_clause_prev[3][49] & ~x[19] & ~x[60] & ~x[61];
			partial_clause[3][50] 	= partial_clause_prev[3][50] & ~x[26];
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & x[62];
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & ~x[22];
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & ~x[51];
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[23] & ~x[54];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & ~x[27];
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & ~x[25];
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & ~x[22];
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & ~x[52];
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & ~x[50];
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & ~x[25];
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & ~x[11];
			partial_clause[4][2] 	= partial_clause_prev[4][2] & ~x[38];
			partial_clause[4][3] 	= partial_clause_prev[4][3] & ~x[11] & ~x[39];
			partial_clause[4][4] 	= partial_clause_prev[4][4] & ~x[10];
			partial_clause[4][5] 	= partial_clause_prev[4][5] & ~x[38];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & ~x[11];
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & ~x[51];
			partial_clause[4][9] 	= partial_clause_prev[4][9] & ~x[10];
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & ~x[10] & ~x[38];
			partial_clause[4][13] 	= partial_clause_prev[4][13] & ~x[38];
			partial_clause[4][14] 	= partial_clause_prev[4][14] & ~x[10] & ~x[38];
			partial_clause[4][15] 	= partial_clause_prev[4][15] & ~x[38];
			partial_clause[4][16] 	= partial_clause_prev[4][16] & ~x[11] & ~x[38];
			partial_clause[4][17] 	= partial_clause_prev[4][17] & ~x[10];
			partial_clause[4][18] 	= partial_clause_prev[4][18] & ~x[10];
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & ~x[38];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & ~x[21] & ~x[38];
			partial_clause[4][23] 	= partial_clause_prev[4][23] & ~x[10];
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & ~x[11];
			partial_clause[4][27] 	= partial_clause_prev[4][27] & ~x[10] & ~x[38];
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & ~x[38];
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[38];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & ~x[11];
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & ~x[38];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & ~x[11];
			partial_clause[4][37] 	= partial_clause_prev[4][37] & ~x[23] & ~x[38] & ~x[48];
			partial_clause[4][38] 	= partial_clause_prev[4][38] & ~x[11] & ~x[38];
			partial_clause[4][39] 	= partial_clause_prev[4][39] & ~x[38];
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & ~x[11];
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & ~x[10];
			partial_clause[4][45] 	= partial_clause_prev[4][45] & ~x[11];
			partial_clause[4][46] 	= partial_clause_prev[4][46] & ~x[39];
			partial_clause[4][47] 	= partial_clause_prev[4][47] & ~x[54];
			partial_clause[4][48] 	= partial_clause_prev[4][48] & ~x[38];
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[11];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & ~x[52];
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & ~x[54];
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & ~x[23];
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & ~x[23];
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & ~x[26];
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & ~x[22];
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & ~x[24];
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & ~x[52];
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & ~x[40] & ~x[41];
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[45];
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & ~x[41] & ~x[42] & ~x[44] & ~x[45] & ~x[46];
			partial_clause[5][7] 	= partial_clause_prev[5][7] & ~x[39] & ~x[40] & ~x[41] & ~x[43] & ~x[44];
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & ~x[42] & ~x[45];
			partial_clause[5][10] 	= partial_clause_prev[5][10] & ~x[41] & ~x[43];
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & ~x[41] & ~x[42] & ~x[45];
			partial_clause[5][16] 	= partial_clause_prev[5][16] & ~x[11] & ~x[12] & ~x[13] & ~x[43] & ~x[44];
			partial_clause[5][17] 	= partial_clause_prev[5][17] & ~x[41] & ~x[45];
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & ~x[40];
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & ~x[42] & ~x[44];
			partial_clause[5][23] 	= partial_clause_prev[5][23] & ~x[42] & ~x[44];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & ~x[25];
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & ~x[39] & ~x[40] & ~x[41] & ~x[43] & ~x[45] & ~x[54];
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & ~x[42] & ~x[43];
			partial_clause[5][31] 	= partial_clause_prev[5][31] & ~x[39] & ~x[41] & ~x[42] & ~x[44];
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & ~x[24] & ~x[40] & ~x[44] & ~x[46];
			partial_clause[5][34] 	= partial_clause_prev[5][34] & ~x[41] & ~x[42] & ~x[44] & ~x[45];
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & ~x[23] & ~x[41];
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & ~x[0] & ~x[41] & ~x[42] & ~x[43];
			partial_clause[5][40] 	= partial_clause_prev[5][40] & ~x[40] & ~x[41] & ~x[42];
			partial_clause[5][41] 	= partial_clause_prev[5][41] & ~x[54];
			partial_clause[5][42] 	= partial_clause_prev[5][42] & ~x[40] & ~x[41];
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & ~x[39] & ~x[40] & ~x[41];
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & ~x[39] & ~x[41];
			partial_clause[5][48] 	= partial_clause_prev[5][48] & ~x[41] & ~x[42];
			partial_clause[5][49] 	= partial_clause_prev[5][49] & ~x[40] & ~x[43] & ~x[44] & ~x[45];
			partial_clause[5][50] 	= partial_clause_prev[5][50] & ~x[19] & ~x[48] & ~x[50];
			partial_clause[5][51] 	= partial_clause_prev[5][51] & ~x[53];
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & ~x[20];
			partial_clause[5][55] 	= partial_clause_prev[5][55] & ~x[47];
			partial_clause[5][56] 	= partial_clause_prev[5][56] & ~x[19] & ~x[48];
			partial_clause[5][57] 	= partial_clause_prev[5][57] & ~x[48];
			partial_clause[5][58] 	= partial_clause_prev[5][58] & ~x[21] & ~x[24];
			partial_clause[5][59] 	= partial_clause_prev[5][59] & ~x[24];
			partial_clause[5][60] 	= partial_clause_prev[5][60] & ~x[19];
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & ~x[19] & ~x[21];
			partial_clause[5][63] 	= partial_clause_prev[5][63] & ~x[18];
			partial_clause[5][64] 	= partial_clause_prev[5][64] & ~x[19] & x[42] & ~x[49];
			partial_clause[5][65] 	= partial_clause_prev[5][65] & ~x[21];
			partial_clause[5][66] 	= partial_clause_prev[5][66] & ~x[20];
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & ~x[48];
			partial_clause[5][69] 	= partial_clause_prev[5][69] & ~x[20] & ~x[21] & x[42] & ~x[48];
			partial_clause[5][70] 	= partial_clause_prev[5][70] & ~x[20] & x[41] & ~x[47];
			partial_clause[5][71] 	= partial_clause_prev[5][71] & ~x[20] & x[43];
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & ~x[47];
			partial_clause[5][74] 	= partial_clause_prev[5][74] & ~x[47];
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & ~x[48];
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & ~x[20];
			partial_clause[5][79] 	= partial_clause_prev[5][79] & ~x[48];
			partial_clause[5][80] 	= partial_clause_prev[5][80] & ~x[19] & ~x[20] & x[42];
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & ~x[19] & ~x[20];
			partial_clause[5][83] 	= partial_clause_prev[5][83] & ~x[21];
			partial_clause[5][84] 	= partial_clause_prev[5][84] & ~x[48];
			partial_clause[5][85] 	= partial_clause_prev[5][85] & ~x[48];
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & x[13] & ~x[21];
			partial_clause[5][88] 	= partial_clause_prev[5][88] & ~x[20];
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & x[42];
			partial_clause[5][91] 	= partial_clause_prev[5][91] & ~x[48] & ~x[50];
			partial_clause[5][92] 	= partial_clause_prev[5][92] & ~x[19];
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & ~x[20];
			partial_clause[5][95] 	= partial_clause_prev[5][95] & ~x[21];
			partial_clause[5][96] 	= partial_clause_prev[5][96] & ~x[49];
			partial_clause[5][97] 	= partial_clause_prev[5][97] & ~x[22];
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & ~x[19] & ~x[48];
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & ~x[13] & ~x[14] & ~x[40];
			partial_clause[6][1] 	= partial_clause_prev[6][1] & ~x[13] & ~x[40];
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & ~x[12] & ~x[14];
			partial_clause[6][4] 	= partial_clause_prev[6][4] & ~x[15] & ~x[40];
			partial_clause[6][5] 	= partial_clause_prev[6][5] & ~x[17];
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & ~x[13];
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & ~x[14] & ~x[40];
			partial_clause[6][10] 	= partial_clause_prev[6][10] & ~x[13];
			partial_clause[6][11] 	= partial_clause_prev[6][11] & ~x[14];
			partial_clause[6][12] 	= partial_clause_prev[6][12] & ~x[14];
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & ~x[13] & ~x[15] & ~x[17] & ~x[40] & ~x[58];
			partial_clause[6][15] 	= partial_clause_prev[6][15] & ~x[12];
			partial_clause[6][16] 	= partial_clause_prev[6][16] & ~x[13] & ~x[16];
			partial_clause[6][17] 	= partial_clause_prev[6][17] & ~x[14] & ~x[40];
			partial_clause[6][18] 	= partial_clause_prev[6][18] & ~x[13] & ~x[15] & ~x[17];
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & ~x[13] & ~x[15] & ~x[19];
			partial_clause[6][21] 	= partial_clause_prev[6][21] & ~x[13];
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & ~x[16] & ~x[41];
			partial_clause[6][25] 	= partial_clause_prev[6][25] & ~x[15] & ~x[41];
			partial_clause[6][26] 	= partial_clause_prev[6][26] & ~x[13] & ~x[15] & ~x[16];
			partial_clause[6][27] 	= partial_clause_prev[6][27] & ~x[49];
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & ~x[13] & ~x[50];
			partial_clause[6][30] 	= partial_clause_prev[6][30] & ~x[40];
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & ~x[15] & ~x[17] & ~x[41] & ~x[55];
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & ~x[40];
			partial_clause[6][35] 	= partial_clause_prev[6][35] & ~x[14];
			partial_clause[6][36] 	= partial_clause_prev[6][36] & ~x[15];
			partial_clause[6][37] 	= partial_clause_prev[6][37] & ~x[40];
			partial_clause[6][38] 	= partial_clause_prev[6][38] & ~x[13];
			partial_clause[6][39] 	= partial_clause_prev[6][39] & ~x[41];
			partial_clause[6][40] 	= partial_clause_prev[6][40] & ~x[13] & ~x[14];
			partial_clause[6][41] 	= partial_clause_prev[6][41] & ~x[13];
			partial_clause[6][42] 	= partial_clause_prev[6][42] & ~x[13] & ~x[16];
			partial_clause[6][43] 	= partial_clause_prev[6][43] & ~x[13] & ~x[16] & ~x[40];
			partial_clause[6][44] 	= partial_clause_prev[6][44] & ~x[40];
			partial_clause[6][45] 	= partial_clause_prev[6][45] & ~x[14] & ~x[16];
			partial_clause[6][46] 	= partial_clause_prev[6][46] & ~x[40];
			partial_clause[6][47] 	= partial_clause_prev[6][47] & ~x[13] & ~x[40] & ~x[41] & ~x[45];
			partial_clause[6][48] 	= partial_clause_prev[6][48] & ~x[15] & ~x[17];
			partial_clause[6][49] 	= partial_clause_prev[6][49] & ~x[54];
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & x[13];
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & ~x[49];
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & x[14];
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & x[16];
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & x[14];
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & ~x[22];
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & ~x[53];
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & ~x[54];
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & ~x[2];
			partial_clause[7][52] 	= partial_clause_prev[7][52] & ~x[23];
			partial_clause[7][53] 	= partial_clause_prev[7][53] & ~x[29];
			partial_clause[7][54] 	= partial_clause_prev[7][54] & ~x[29];
			partial_clause[7][55] 	= partial_clause_prev[7][55] & ~x[30] & ~x[57];
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & ~x[56];
			partial_clause[7][60] 	= partial_clause_prev[7][60] & ~x[57];
			partial_clause[7][61] 	= partial_clause_prev[7][61] & ~x[52];
			partial_clause[7][62] 	= partial_clause_prev[7][62] & ~x[28];
			partial_clause[7][63] 	= partial_clause_prev[7][63] & ~x[55];
			partial_clause[7][64] 	= partial_clause_prev[7][64] & ~x[2] & ~x[27];
			partial_clause[7][65] 	= partial_clause_prev[7][65] & ~x[3];
			partial_clause[7][66] 	= partial_clause_prev[7][66] & ~x[2];
			partial_clause[7][67] 	= partial_clause_prev[7][67] & ~x[56];
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & ~x[1] & ~x[28];
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & ~x[2];
			partial_clause[7][73] 	= partial_clause_prev[7][73] & ~x[41] & ~x[56];
			partial_clause[7][74] 	= partial_clause_prev[7][74] & ~x[30];
			partial_clause[7][75] 	= partial_clause_prev[7][75] & ~x[28];
			partial_clause[7][76] 	= partial_clause_prev[7][76] & ~x[30];
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & ~x[56];
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & ~x[28];
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & ~x[30];
			partial_clause[7][85] 	= partial_clause_prev[7][85] & ~x[1];
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & ~x[2];
			partial_clause[7][89] 	= partial_clause_prev[7][89] & ~x[57];
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & ~x[3] & ~x[28];
			partial_clause[7][93] 	= partial_clause_prev[7][93] & ~x[29];
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & ~x[31];
			partial_clause[7][96] 	= partial_clause_prev[7][96] & ~x[1];
			partial_clause[7][97] 	= partial_clause_prev[7][97] & ~x[28];
			partial_clause[7][98] 	= partial_clause_prev[7][98] & ~x[1] & ~x[57];
			partial_clause[7][99] 	= partial_clause_prev[7][99] & ~x[28];
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & ~x[55] & x[63];
			partial_clause[8][6] 	= partial_clause_prev[8][6] & ~x[55];
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & ~x[0];
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & ~x[28];
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & ~x[11] & ~x[25];
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & x[35];
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & ~x[55];
			partial_clause[8][27] 	= partial_clause_prev[8][27] & ~x[1];
			partial_clause[8][28] 	= partial_clause_prev[8][28] & ~x[27];
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & ~x[1];
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & ~x[11];
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & ~x[38];
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & ~x[49];
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & ~x[20];
			partial_clause[8][55] 	= partial_clause_prev[8][55] & ~x[20] & ~x[23];
			partial_clause[8][56] 	= partial_clause_prev[8][56] & ~x[18] & ~x[47];
			partial_clause[8][57] 	= partial_clause_prev[8][57] & ~x[20];
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & ~x[20] & ~x[50];
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & ~x[18];
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & ~x[20];
			partial_clause[8][64] 	= partial_clause_prev[8][64] & ~x[20];
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & ~x[20] & ~x[49];
			partial_clause[8][67] 	= partial_clause_prev[8][67] & ~x[21];
			partial_clause[8][68] 	= partial_clause_prev[8][68] & ~x[49];
			partial_clause[8][69] 	= partial_clause_prev[8][69] & ~x[47];
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & ~x[18] & ~x[19];
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & ~x[49];
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & ~x[47];
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & ~x[20];
			partial_clause[8][80] 	= partial_clause_prev[8][80] & ~x[20] & ~x[23];
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & ~x[46] & ~x[47];
			partial_clause[8][83] 	= partial_clause_prev[8][83] & ~x[19];
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & ~x[20];
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & ~x[20];
			partial_clause[8][89] 	= partial_clause_prev[8][89] & ~x[48];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & ~x[47] & ~x[52];
			partial_clause[8][92] 	= partial_clause_prev[8][92] & ~x[0] & ~x[20] & ~x[47];
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & ~x[17] & ~x[29] & ~x[32] & ~x[33] & ~x[45];
			partial_clause[8][95] 	= partial_clause_prev[8][95] & ~x[49];
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & ~x[20];
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & ~x[53];
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & ~x[2];
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & ~x[2];
			partial_clause[9][6] 	= partial_clause_prev[9][6] & ~x[27];
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & ~x[3];
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & ~x[2];
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & ~x[2];
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & ~x[24];
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & ~x[28];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & ~x[1];
			partial_clause[9][42] 	= partial_clause_prev[9][42] & ~x[0];
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & ~x[29];
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & ~x[2];
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & ~x[50];
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & ~x[52] & ~x[54];
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & ~x[27];
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & ~x[21];
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & ~x[33] & ~x[61] & ~x[62];
			partial_clause[9][67] 	= partial_clause_prev[9][67] & ~x[54];
			partial_clause[9][68] 	= partial_clause_prev[9][68] & ~x[56];
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & ~x[62];
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
		end
	end
endmodule


module HCB_5 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & ~x[19];
			partial_clause[0][2] 	= partial_clause_prev[0][2] & ~x[60];
			partial_clause[0][3] 	= partial_clause_prev[0][3] & ~x[60];
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & ~x[17] & ~x[32];
			partial_clause[0][6] 	= partial_clause_prev[0][6] & ~x[31];
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & ~x[30];
			partial_clause[0][9] 	= partial_clause_prev[0][9] & ~x[32];
			partial_clause[0][10] 	= partial_clause_prev[0][10] & ~x[31];
			partial_clause[0][11] 	= partial_clause_prev[0][11] & ~x[31] & ~x[59];
			partial_clause[0][12] 	= partial_clause_prev[0][12] & ~x[31] & ~x[59];
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & ~x[59];
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & ~x[58] & ~x[61];
			partial_clause[0][17] 	= partial_clause_prev[0][17] & ~x[31] & ~x[32] & ~x[58];
			partial_clause[0][18] 	= partial_clause_prev[0][18] & ~x[43] & ~x[60];
			partial_clause[0][19] 	= partial_clause_prev[0][19] & ~x[61];
			partial_clause[0][20] 	= partial_clause_prev[0][20] & ~x[32] & ~x[59];
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & ~x[32] & ~x[60];
			partial_clause[0][23] 	= partial_clause_prev[0][23] & ~x[60];
			partial_clause[0][24] 	= partial_clause_prev[0][24] & ~x[32] & ~x[33];
			partial_clause[0][25] 	= partial_clause_prev[0][25] & ~x[32];
			partial_clause[0][26] 	= partial_clause_prev[0][26] & ~x[57] & ~x[60];
			partial_clause[0][27] 	= partial_clause_prev[0][27] & ~x[4];
			partial_clause[0][28] 	= partial_clause_prev[0][28] & ~x[61];
			partial_clause[0][29] 	= partial_clause_prev[0][29] & ~x[60];
			partial_clause[0][30] 	= partial_clause_prev[0][30] & ~x[60];
			partial_clause[0][31] 	= partial_clause_prev[0][31] & ~x[58];
			partial_clause[0][32] 	= partial_clause_prev[0][32] & ~x[31];
			partial_clause[0][33] 	= partial_clause_prev[0][33] & ~x[31];
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & ~x[59];
			partial_clause[0][36] 	= partial_clause_prev[0][36] & ~x[32] & ~x[59];
			partial_clause[0][37] 	= partial_clause_prev[0][37] & ~x[31];
			partial_clause[0][38] 	= partial_clause_prev[0][38] & ~x[32];
			partial_clause[0][39] 	= partial_clause_prev[0][39] & ~x[31];
			partial_clause[0][40] 	= partial_clause_prev[0][40] & ~x[32];
			partial_clause[0][41] 	= partial_clause_prev[0][41] & ~x[58];
			partial_clause[0][42] 	= partial_clause_prev[0][42] & ~x[31] & ~x[60];
			partial_clause[0][43] 	= partial_clause_prev[0][43] & ~x[32] & ~x[60];
			partial_clause[0][44] 	= partial_clause_prev[0][44] & ~x[32];
			partial_clause[0][45] 	= partial_clause_prev[0][45] & ~x[31] & ~x[45];
			partial_clause[0][46] 	= partial_clause_prev[0][46] & ~x[58] & ~x[61];
			partial_clause[0][47] 	= partial_clause_prev[0][47] & ~x[59] & ~x[61];
			partial_clause[0][48] 	= partial_clause_prev[0][48] & ~x[32];
			partial_clause[0][49] 	= partial_clause_prev[0][49] & ~x[59];
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & ~x[46];
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & ~x[39];
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & ~x[11] & ~x[44];
			partial_clause[0][58] 	= partial_clause_prev[0][58] & ~x[39];
			partial_clause[0][59] 	= partial_clause_prev[0][59] & ~x[18];
			partial_clause[0][60] 	= partial_clause_prev[0][60] & ~x[19];
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & ~x[11];
			partial_clause[0][63] 	= partial_clause_prev[0][63] & ~x[11] & ~x[36] & ~x[44];
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & ~x[40];
			partial_clause[0][66] 	= partial_clause_prev[0][66] & ~x[39];
			partial_clause[0][67] 	= partial_clause_prev[0][67] & ~x[18] & ~x[46];
			partial_clause[0][68] 	= partial_clause_prev[0][68] & ~x[41];
			partial_clause[0][69] 	= partial_clause_prev[0][69] & ~x[43];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & ~x[36];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & ~x[39];
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & ~x[15];
			partial_clause[0][74] 	= partial_clause_prev[0][74] & ~x[11];
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & ~x[38];
			partial_clause[0][78] 	= partial_clause_prev[0][78] & ~x[11] & x[59];
			partial_clause[0][79] 	= partial_clause_prev[0][79] & ~x[40] & ~x[41];
			partial_clause[0][80] 	= partial_clause_prev[0][80] & ~x[11];
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & ~x[40];
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & ~x[39] & x[60];
			partial_clause[0][86] 	= partial_clause_prev[0][86] & ~x[44];
			partial_clause[0][87] 	= partial_clause_prev[0][87] & ~x[10] & ~x[14];
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & ~x[11];
			partial_clause[0][90] 	= partial_clause_prev[0][90] & ~x[38] & ~x[40];
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & ~x[38];
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & ~x[35] & ~x[37];
			partial_clause[0][96] 	= partial_clause_prev[0][96] & ~x[38];
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & ~x[38];
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[23] & ~x[27];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & ~x[8] & ~x[35];
			partial_clause[1][2] 	= partial_clause_prev[1][2] & x[58];
			partial_clause[1][3] 	= partial_clause_prev[1][3] & ~x[34];
			partial_clause[1][4] 	= partial_clause_prev[1][4] & ~x[26];
			partial_clause[1][5] 	= partial_clause_prev[1][5] & ~x[8] & ~x[54];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & ~x[22];
			partial_clause[1][7] 	= partial_clause_prev[1][7] & x[30] & ~x[55];
			partial_clause[1][8] 	= partial_clause_prev[1][8] & ~x[27];
			partial_clause[1][9] 	= partial_clause_prev[1][9] & ~x[7] & ~x[26];
			partial_clause[1][10] 	= partial_clause_prev[1][10] & ~x[9];
			partial_clause[1][11] 	= partial_clause_prev[1][11] & ~x[8] & ~x[55] & x[58];
			partial_clause[1][12] 	= partial_clause_prev[1][12] & ~x[26];
			partial_clause[1][13] 	= partial_clause_prev[1][13] & x[58];
			partial_clause[1][14] 	= partial_clause_prev[1][14] & x[30] & ~x[35] & ~x[54];
			partial_clause[1][15] 	= partial_clause_prev[1][15] & x[30];
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & ~x[27] & x[58];
			partial_clause[1][18] 	= partial_clause_prev[1][18] & x[30] & ~x[54];
			partial_clause[1][19] 	= partial_clause_prev[1][19] & x[58];
			partial_clause[1][20] 	= partial_clause_prev[1][20] & x[30] & ~x[54] & ~x[62];
			partial_clause[1][21] 	= partial_clause_prev[1][21] & ~x[9] & ~x[35] & ~x[62];
			partial_clause[1][22] 	= partial_clause_prev[1][22] & ~x[54];
			partial_clause[1][23] 	= partial_clause_prev[1][23] & ~x[8] & ~x[25] & x[30] & ~x[55];
			partial_clause[1][24] 	= partial_clause_prev[1][24] & ~x[35] & ~x[52];
			partial_clause[1][25] 	= partial_clause_prev[1][25] & ~x[55] & x[58] & ~x[62];
			partial_clause[1][26] 	= partial_clause_prev[1][26] & x[30];
			partial_clause[1][27] 	= partial_clause_prev[1][27] & ~x[53] & x[58];
			partial_clause[1][28] 	= partial_clause_prev[1][28] & x[58];
			partial_clause[1][29] 	= partial_clause_prev[1][29] & ~x[27];
			partial_clause[1][30] 	= partial_clause_prev[1][30] & x[30] & ~x[55];
			partial_clause[1][31] 	= partial_clause_prev[1][31] & ~x[27];
			partial_clause[1][32] 	= partial_clause_prev[1][32] & ~x[25] & ~x[26] & x[58];
			partial_clause[1][33] 	= partial_clause_prev[1][33] & ~x[23];
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & ~x[55];
			partial_clause[1][36] 	= partial_clause_prev[1][36] & ~x[35] & ~x[55];
			partial_clause[1][37] 	= partial_clause_prev[1][37] & x[30];
			partial_clause[1][38] 	= partial_clause_prev[1][38] & ~x[27] & ~x[55];
			partial_clause[1][39] 	= partial_clause_prev[1][39] & ~x[26] & x[58];
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & ~x[55] & x[58];
			partial_clause[1][42] 	= partial_clause_prev[1][42] & x[58];
			partial_clause[1][43] 	= partial_clause_prev[1][43] & x[58];
			partial_clause[1][44] 	= partial_clause_prev[1][44] & ~x[55];
			partial_clause[1][45] 	= partial_clause_prev[1][45] & ~x[62];
			partial_clause[1][46] 	= partial_clause_prev[1][46] & ~x[27] & ~x[61];
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & ~x[33] & ~x[54];
			partial_clause[1][49] 	= partial_clause_prev[1][49] & ~x[7] & ~x[55];
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & ~x[30];
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & x[34];
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & ~x[45];
			partial_clause[1][56] 	= partial_clause_prev[1][56] & ~x[16] & ~x[30] & ~x[31];
			partial_clause[1][57] 	= partial_clause_prev[1][57] & x[55];
			partial_clause[1][58] 	= partial_clause_prev[1][58] & 1'b1;
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & ~x[58];
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & ~x[3] & ~x[18] & ~x[44] & ~x[46];
			partial_clause[1][64] 	= partial_clause_prev[1][64] & ~x[30];
			partial_clause[1][65] 	= partial_clause_prev[1][65] & ~x[3];
			partial_clause[1][66] 	= partial_clause_prev[1][66] & ~x[30];
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & x[27] & ~x[43];
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & x[25];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & ~x[45];
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & ~x[30];
			partial_clause[1][80] 	= partial_clause_prev[1][80] & ~x[13] & ~x[45];
			partial_clause[1][81] 	= partial_clause_prev[1][81] & ~x[2] & ~x[3] & ~x[17];
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & ~x[46];
			partial_clause[1][87] 	= partial_clause_prev[1][87] & ~x[17];
			partial_clause[1][88] 	= partial_clause_prev[1][88] & ~x[2] & ~x[3] & ~x[45];
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & ~x[16] & x[55];
			partial_clause[1][91] 	= partial_clause_prev[1][91] & ~x[18] & ~x[47];
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & x[26];
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & ~x[15] & x[34];
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & ~x[51] & ~x[52];
			partial_clause[2][1] 	= partial_clause_prev[2][1] & ~x[1] & ~x[27] & ~x[29] & ~x[30] & ~x[43] & ~x[51];
			partial_clause[2][2] 	= partial_clause_prev[2][2] & ~x[0] & ~x[1] & ~x[2] & ~x[24] & ~x[26] & ~x[50];
			partial_clause[2][3] 	= partial_clause_prev[2][3] & ~x[1] & ~x[13] & ~x[27];
			partial_clause[2][4] 	= partial_clause_prev[2][4] & ~x[50] & ~x[52];
			partial_clause[2][5] 	= partial_clause_prev[2][5] & ~x[0] & ~x[2] & ~x[24] & ~x[26];
			partial_clause[2][6] 	= partial_clause_prev[2][6] & ~x[0] & ~x[24];
			partial_clause[2][7] 	= partial_clause_prev[2][7] & ~x[0];
			partial_clause[2][8] 	= partial_clause_prev[2][8] & ~x[0] & ~x[1] & ~x[24] & ~x[27] & ~x[52];
			partial_clause[2][9] 	= partial_clause_prev[2][9] & ~x[26] & ~x[27] & ~x[50];
			partial_clause[2][10] 	= partial_clause_prev[2][10] & ~x[2] & ~x[23];
			partial_clause[2][11] 	= partial_clause_prev[2][11] & ~x[0] & ~x[23] & ~x[26] & ~x[29];
			partial_clause[2][12] 	= partial_clause_prev[2][12] & ~x[1] & ~x[25] & ~x[26] & ~x[50];
			partial_clause[2][13] 	= partial_clause_prev[2][13] & ~x[23] & ~x[25];
			partial_clause[2][14] 	= partial_clause_prev[2][14] & ~x[26] & ~x[52];
			partial_clause[2][15] 	= partial_clause_prev[2][15] & ~x[1] & ~x[13] & ~x[23] & ~x[25] & ~x[26];
			partial_clause[2][16] 	= partial_clause_prev[2][16] & ~x[24] & ~x[25] & ~x[26] & ~x[30];
			partial_clause[2][17] 	= partial_clause_prev[2][17] & ~x[1] & ~x[23];
			partial_clause[2][18] 	= partial_clause_prev[2][18] & ~x[1] & ~x[27] & ~x[51];
			partial_clause[2][19] 	= partial_clause_prev[2][19] & ~x[1] & ~x[22] & ~x[26] & ~x[27] & ~x[51];
			partial_clause[2][20] 	= partial_clause_prev[2][20] & ~x[22] & ~x[25] & ~x[27] & ~x[30] & ~x[52];
			partial_clause[2][21] 	= partial_clause_prev[2][21] & ~x[23] & ~x[24] & ~x[26] & ~x[27] & ~x[28];
			partial_clause[2][22] 	= partial_clause_prev[2][22] & ~x[27] & ~x[28] & ~x[49] & ~x[50] & ~x[51];
			partial_clause[2][23] 	= partial_clause_prev[2][23] & ~x[2] & ~x[23] & ~x[25] & ~x[26] & ~x[52];
			partial_clause[2][24] 	= partial_clause_prev[2][24] & ~x[14] & ~x[23] & ~x[42];
			partial_clause[2][25] 	= partial_clause_prev[2][25] & ~x[25] & ~x[27] & ~x[28];
			partial_clause[2][26] 	= partial_clause_prev[2][26] & ~x[26] & ~x[27] & ~x[51];
			partial_clause[2][27] 	= partial_clause_prev[2][27] & ~x[0] & ~x[1] & ~x[2] & ~x[23];
			partial_clause[2][28] 	= partial_clause_prev[2][28] & ~x[1] & ~x[24];
			partial_clause[2][29] 	= partial_clause_prev[2][29] & ~x[2] & ~x[23] & ~x[27] & ~x[49] & ~x[53];
			partial_clause[2][30] 	= partial_clause_prev[2][30] & ~x[1] & ~x[23] & ~x[26] & ~x[52];
			partial_clause[2][31] 	= partial_clause_prev[2][31] & ~x[1] & ~x[22] & ~x[28];
			partial_clause[2][32] 	= partial_clause_prev[2][32] & ~x[1] & ~x[27] & ~x[52];
			partial_clause[2][33] 	= partial_clause_prev[2][33] & ~x[13] & ~x[25] & ~x[27];
			partial_clause[2][34] 	= partial_clause_prev[2][34] & ~x[0] & ~x[2] & ~x[25] & ~x[27];
			partial_clause[2][35] 	= partial_clause_prev[2][35] & ~x[1] & ~x[24] & ~x[28] & ~x[51];
			partial_clause[2][36] 	= partial_clause_prev[2][36] & ~x[23] & ~x[26] & ~x[29];
			partial_clause[2][37] 	= partial_clause_prev[2][37] & ~x[1] & ~x[22] & ~x[28] & ~x[39];
			partial_clause[2][38] 	= partial_clause_prev[2][38] & ~x[24] & ~x[29] & ~x[50] & ~x[54];
			partial_clause[2][39] 	= partial_clause_prev[2][39] & ~x[0] & ~x[2] & ~x[26] & ~x[52];
			partial_clause[2][40] 	= partial_clause_prev[2][40] & ~x[22] & ~x[25];
			partial_clause[2][41] 	= partial_clause_prev[2][41] & ~x[0] & ~x[27] & ~x[48] & ~x[51] & ~x[52];
			partial_clause[2][42] 	= partial_clause_prev[2][42] & ~x[0] & ~x[1];
			partial_clause[2][43] 	= partial_clause_prev[2][43] & ~x[24] & ~x[26] & ~x[53];
			partial_clause[2][44] 	= partial_clause_prev[2][44] & ~x[0] & ~x[24] & ~x[26];
			partial_clause[2][45] 	= partial_clause_prev[2][45] & ~x[1] & ~x[22] & ~x[24];
			partial_clause[2][46] 	= partial_clause_prev[2][46] & ~x[23] & ~x[27] & ~x[29];
			partial_clause[2][47] 	= partial_clause_prev[2][47] & ~x[0] & ~x[23] & ~x[26];
			partial_clause[2][48] 	= partial_clause_prev[2][48] & ~x[0] & ~x[24] & ~x[50];
			partial_clause[2][49] 	= partial_clause_prev[2][49] & ~x[0] & ~x[1] & ~x[2] & ~x[24] & ~x[25];
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & x[53];
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & ~x[41];
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & ~x[15];
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & x[27];
			partial_clause[2][65] 	= partial_clause_prev[2][65] & ~x[41];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & ~x[21] & x[27];
			partial_clause[2][68] 	= partial_clause_prev[2][68] & ~x[19] & x[27];
			partial_clause[2][69] 	= partial_clause_prev[2][69] & x[26];
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & x[26] & ~x[42];
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & ~x[47];
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & ~x[41];
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & x[27];
			partial_clause[2][80] 	= partial_clause_prev[2][80] & ~x[13];
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & x[25] & ~x[42];
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & x[54];
			partial_clause[2][89] 	= partial_clause_prev[2][89] & ~x[44] & x[53];
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & x[26];
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & x[53];
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & ~x[23] & x[30];
			partial_clause[3][2] 	= partial_clause_prev[3][2] & x[30];
			partial_clause[3][3] 	= partial_clause_prev[3][3] & x[30];
			partial_clause[3][4] 	= partial_clause_prev[3][4] & x[30] & ~x[40];
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & ~x[37];
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & ~x[11];
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & ~x[49];
			partial_clause[3][13] 	= partial_clause_prev[3][13] & ~x[15];
			partial_clause[3][14] 	= partial_clause_prev[3][14] & ~x[38];
			partial_clause[3][15] 	= partial_clause_prev[3][15] & ~x[50];
			partial_clause[3][16] 	= partial_clause_prev[3][16] & ~x[14] & ~x[51] & x[57];
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & ~x[37];
			partial_clause[3][21] 	= partial_clause_prev[3][21] & ~x[23];
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & x[31] & ~x[51];
			partial_clause[3][24] 	= partial_clause_prev[3][24] & ~x[22];
			partial_clause[3][25] 	= partial_clause_prev[3][25] & ~x[10];
			partial_clause[3][26] 	= partial_clause_prev[3][26] & x[30];
			partial_clause[3][27] 	= partial_clause_prev[3][27] & ~x[23];
			partial_clause[3][28] 	= partial_clause_prev[3][28] & ~x[23];
			partial_clause[3][29] 	= partial_clause_prev[3][29] & ~x[23];
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & x[30];
			partial_clause[3][32] 	= partial_clause_prev[3][32] & ~x[39];
			partial_clause[3][33] 	= partial_clause_prev[3][33] & ~x[10];
			partial_clause[3][34] 	= partial_clause_prev[3][34] & ~x[23] & ~x[40];
			partial_clause[3][35] 	= partial_clause_prev[3][35] & ~x[24] & x[58];
			partial_clause[3][36] 	= partial_clause_prev[3][36] & ~x[22] & x[31];
			partial_clause[3][37] 	= partial_clause_prev[3][37] & ~x[22];
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & x[57];
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & x[30] & x[31];
			partial_clause[3][46] 	= partial_clause_prev[3][46] & ~x[39];
			partial_clause[3][47] 	= partial_clause_prev[3][47] & ~x[22];
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & ~x[29] & ~x[57];
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & ~x[30] & ~x[31] & ~x[46];
			partial_clause[3][54] 	= partial_clause_prev[3][54] & ~x[56];
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & ~x[2] & ~x[30];
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & ~x[3] & ~x[31];
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & ~x[30] & ~x[58];
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[30];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & ~x[29] & ~x[30];
			partial_clause[3][67] 	= partial_clause_prev[3][67] & ~x[30] & ~x[58];
			partial_clause[3][68] 	= partial_clause_prev[3][68] & ~x[4];
			partial_clause[3][69] 	= partial_clause_prev[3][69] & ~x[3] & ~x[58];
			partial_clause[3][70] 	= partial_clause_prev[3][70] & ~x[3] & ~x[16];
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & ~x[30] & ~x[57];
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & ~x[30];
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & ~x[30];
			partial_clause[3][79] 	= partial_clause_prev[3][79] & ~x[42];
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & ~x[43] & ~x[58];
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & ~x[31];
			partial_clause[3][86] 	= partial_clause_prev[3][86] & ~x[4];
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & ~x[19];
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & ~x[2] & ~x[14] & ~x[30];
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & ~x[17];
			partial_clause[3][95] 	= partial_clause_prev[3][95] & ~x[2] & ~x[30];
			partial_clause[3][96] 	= partial_clause_prev[3][96] & ~x[3] & ~x[31];
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & ~x[3];
			partial_clause[4][2] 	= partial_clause_prev[4][2] & ~x[2] & ~x[43];
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & ~x[30];
			partial_clause[4][11] 	= partial_clause_prev[4][11] & ~x[2];
			partial_clause[4][12] 	= partial_clause_prev[4][12] & ~x[13];
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & ~x[2];
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & ~x[2];
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & ~x[2];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & ~x[2];
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & ~x[2];
			partial_clause[4][31] 	= partial_clause_prev[4][31] & ~x[2];
			partial_clause[4][32] 	= partial_clause_prev[4][32] & 1'b1;
			partial_clause[4][33] 	= partial_clause_prev[4][33] & ~x[2];
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & ~x[2];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & ~x[2];
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & ~x[2];
			partial_clause[4][41] 	= partial_clause_prev[4][41] & ~x[2];
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & ~x[47];
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & 1'b1;
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & ~x[53];
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & ~x[44] & ~x[52];
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & ~x[52] & ~x[54];
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & ~x[45];
			partial_clause[4][69] 	= partial_clause_prev[4][69] & ~x[48];
			partial_clause[4][70] 	= partial_clause_prev[4][70] & ~x[20];
			partial_clause[4][71] 	= partial_clause_prev[4][71] & ~x[51] & ~x[53];
			partial_clause[4][72] 	= partial_clause_prev[4][72] & ~x[13];
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & ~x[54];
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & ~x[42];
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & ~x[19];
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & ~x[41] & ~x[42] & ~x[53];
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & ~x[15];
			partial_clause[4][95] 	= partial_clause_prev[4][95] & ~x[19];
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & ~x[5] & ~x[6] & ~x[17];
			partial_clause[5][1] 	= partial_clause_prev[5][1] & ~x[7];
			partial_clause[5][2] 	= partial_clause_prev[5][2] & ~x[4] & ~x[35];
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & ~x[31] & ~x[33] & ~x[45] & ~x[63];
			partial_clause[5][5] 	= partial_clause_prev[5][5] & ~x[3] & ~x[5] & ~x[7] & ~x[8] & ~x[10];
			partial_clause[5][6] 	= partial_clause_prev[5][6] & ~x[9];
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & ~x[5] & ~x[6] & ~x[8];
			partial_clause[5][9] 	= partial_clause_prev[5][9] & ~x[7] & ~x[8] & ~x[37];
			partial_clause[5][10] 	= partial_clause_prev[5][10] & ~x[9];
			partial_clause[5][11] 	= partial_clause_prev[5][11] & ~x[3] & ~x[8] & ~x[34] & ~x[39];
			partial_clause[5][12] 	= partial_clause_prev[5][12] & ~x[33] & ~x[34] & x[55];
			partial_clause[5][13] 	= partial_clause_prev[5][13] & ~x[3] & ~x[35] & ~x[37];
			partial_clause[5][14] 	= partial_clause_prev[5][14] & ~x[4] & ~x[5] & ~x[6] & ~x[8] & ~x[9];
			partial_clause[5][15] 	= partial_clause_prev[5][15] & ~x[7] & ~x[10];
			partial_clause[5][16] 	= partial_clause_prev[5][16] & ~x[9];
			partial_clause[5][17] 	= partial_clause_prev[5][17] & ~x[10] & ~x[11];
			partial_clause[5][18] 	= partial_clause_prev[5][18] & ~x[6] & ~x[36] & ~x[45] & x[54];
			partial_clause[5][19] 	= partial_clause_prev[5][19] & ~x[6];
			partial_clause[5][20] 	= partial_clause_prev[5][20] & ~x[4] & ~x[5] & ~x[7] & ~x[39];
			partial_clause[5][21] 	= partial_clause_prev[5][21] & ~x[35] & ~x[36] & ~x[38];
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & ~x[9];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & ~x[5] & ~x[7] & ~x[38];
			partial_clause[5][25] 	= partial_clause_prev[5][25] & ~x[4] & ~x[6] & ~x[7] & ~x[36] & x[55];
			partial_clause[5][26] 	= partial_clause_prev[5][26] & ~x[6] & ~x[8] & ~x[9] & ~x[37];
			partial_clause[5][27] 	= partial_clause_prev[5][27] & ~x[7] & x[27] & ~x[42];
			partial_clause[5][28] 	= partial_clause_prev[5][28] & ~x[7];
			partial_clause[5][29] 	= partial_clause_prev[5][29] & ~x[3] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[36] & ~x[39];
			partial_clause[5][30] 	= partial_clause_prev[5][30] & ~x[8];
			partial_clause[5][31] 	= partial_clause_prev[5][31] & ~x[9];
			partial_clause[5][32] 	= partial_clause_prev[5][32] & ~x[5] & ~x[6] & ~x[7] & ~x[39] & x[55];
			partial_clause[5][33] 	= partial_clause_prev[5][33] & ~x[7] & ~x[37];
			partial_clause[5][34] 	= partial_clause_prev[5][34] & ~x[11];
			partial_clause[5][35] 	= partial_clause_prev[5][35] & ~x[4] & ~x[6] & ~x[8] & x[55];
			partial_clause[5][36] 	= partial_clause_prev[5][36] & ~x[8] & ~x[38];
			partial_clause[5][37] 	= partial_clause_prev[5][37] & ~x[4] & ~x[7] & ~x[9] & ~x[10] & ~x[35];
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & ~x[9] & ~x[39];
			partial_clause[5][40] 	= partial_clause_prev[5][40] & ~x[9];
			partial_clause[5][41] 	= partial_clause_prev[5][41] & ~x[6] & ~x[7] & ~x[9] & x[26] & ~x[45];
			partial_clause[5][42] 	= partial_clause_prev[5][42] & ~x[7] & ~x[9];
			partial_clause[5][43] 	= partial_clause_prev[5][43] & ~x[8] & ~x[36] & ~x[38];
			partial_clause[5][44] 	= partial_clause_prev[5][44] & ~x[31] & ~x[62];
			partial_clause[5][45] 	= partial_clause_prev[5][45] & ~x[8] & ~x[16] & ~x[37];
			partial_clause[5][46] 	= partial_clause_prev[5][46] & ~x[6] & x[27] & ~x[36] & ~x[41];
			partial_clause[5][47] 	= partial_clause_prev[5][47] & ~x[6] & ~x[9] & ~x[10];
			partial_clause[5][48] 	= partial_clause_prev[5][48] & ~x[7] & ~x[37] & ~x[38];
			partial_clause[5][49] 	= partial_clause_prev[5][49] & ~x[11];
			partial_clause[5][50] 	= partial_clause_prev[5][50] & ~x[44];
			partial_clause[5][51] 	= partial_clause_prev[5][51] & x[62];
			partial_clause[5][52] 	= partial_clause_prev[5][52] & ~x[27];
			partial_clause[5][53] 	= partial_clause_prev[5][53] & ~x[2] & x[6];
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & ~x[16] & ~x[27];
			partial_clause[5][57] 	= partial_clause_prev[5][57] & ~x[26];
			partial_clause[5][58] 	= partial_clause_prev[5][58] & ~x[28];
			partial_clause[5][59] 	= partial_clause_prev[5][59] & x[6] & ~x[44];
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & x[32];
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & ~x[41];
			partial_clause[5][65] 	= partial_clause_prev[5][65] & ~x[28] & ~x[46] & ~x[56];
			partial_clause[5][66] 	= partial_clause_prev[5][66] & ~x[27];
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & ~x[0] & ~x[55];
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & ~x[28] & ~x[55];
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & x[61];
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & ~x[13];
			partial_clause[5][80] 	= partial_clause_prev[5][80] & ~x[12];
			partial_clause[5][81] 	= partial_clause_prev[5][81] & ~x[3] & x[35];
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & ~x[27];
			partial_clause[5][84] 	= partial_clause_prev[5][84] & ~x[12];
			partial_clause[5][85] 	= partial_clause_prev[5][85] & ~x[27] & ~x[55];
			partial_clause[5][86] 	= partial_clause_prev[5][86] & ~x[0] & ~x[55];
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & ~x[12] & ~x[13];
			partial_clause[5][89] 	= partial_clause_prev[5][89] & ~x[0] & ~x[55];
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & x[5];
			partial_clause[5][92] 	= partial_clause_prev[5][92] & ~x[26];
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & ~x[0] & ~x[27];
			partial_clause[5][95] 	= partial_clause_prev[5][95] & ~x[30] & x[34];
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & x[33];
			partial_clause[5][98] 	= partial_clause_prev[5][98] & ~x[27];
			partial_clause[5][99] 	= partial_clause_prev[5][99] & ~x[28];
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & ~x[14];
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & ~x[20] & ~x[21];
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & ~x[41];
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & ~x[47];
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & ~x[18];
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & ~x[3];
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & ~x[17];
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & ~x[44];
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & x[55];
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & ~x[47];
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & ~x[18];
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & ~x[47];
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & ~x[45];
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & ~x[14];
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & ~x[57];
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & ~x[17] & ~x[57];
			partial_clause[7][3] 	= partial_clause_prev[7][3] & ~x[57];
			partial_clause[7][4] 	= partial_clause_prev[7][4] & ~x[58];
			partial_clause[7][5] 	= partial_clause_prev[7][5] & ~x[57];
			partial_clause[7][6] 	= partial_clause_prev[7][6] & ~x[57];
			partial_clause[7][7] 	= partial_clause_prev[7][7] & ~x[13];
			partial_clause[7][8] 	= partial_clause_prev[7][8] & ~x[58];
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & ~x[30];
			partial_clause[7][11] 	= partial_clause_prev[7][11] & ~x[57];
			partial_clause[7][12] 	= partial_clause_prev[7][12] & ~x[58];
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & ~x[58];
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & ~x[57];
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & ~x[57];
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & ~x[57];
			partial_clause[7][21] 	= partial_clause_prev[7][21] & ~x[58];
			partial_clause[7][22] 	= partial_clause_prev[7][22] & ~x[57];
			partial_clause[7][23] 	= partial_clause_prev[7][23] & ~x[57];
			partial_clause[7][24] 	= partial_clause_prev[7][24] & ~x[57];
			partial_clause[7][25] 	= partial_clause_prev[7][25] & ~x[30];
			partial_clause[7][26] 	= partial_clause_prev[7][26] & ~x[57] & ~x[58];
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & ~x[57];
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & ~x[57];
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & ~x[57];
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & ~x[57];
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & ~x[57] & ~x[58];
			partial_clause[7][40] 	= partial_clause_prev[7][40] & ~x[57];
			partial_clause[7][41] 	= partial_clause_prev[7][41] & ~x[57];
			partial_clause[7][42] 	= partial_clause_prev[7][42] & ~x[57] & ~x[58];
			partial_clause[7][43] 	= partial_clause_prev[7][43] & ~x[57];
			partial_clause[7][44] 	= partial_clause_prev[7][44] & ~x[57];
			partial_clause[7][45] 	= partial_clause_prev[7][45] & ~x[57];
			partial_clause[7][46] 	= partial_clause_prev[7][46] & ~x[57];
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & ~x[58];
			partial_clause[7][49] 	= partial_clause_prev[7][49] & ~x[58];
			partial_clause[7][50] 	= partial_clause_prev[7][50] & ~x[14];
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & ~x[18];
			partial_clause[7][54] 	= partial_clause_prev[7][54] & ~x[14];
			partial_clause[7][55] 	= partial_clause_prev[7][55] & ~x[48];
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & ~x[20];
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & ~x[42];
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & x[57];
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & ~x[19] & ~x[20];
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & ~x[46];
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & ~x[20] & x[57];
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & x[58];
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & ~x[20];
			partial_clause[7][86] 	= partial_clause_prev[7][86] & ~x[21] & x[56];
			partial_clause[7][87] 	= partial_clause_prev[7][87] & ~x[21];
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & ~x[20] & x[55];
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & ~x[20];
			partial_clause[7][97] 	= partial_clause_prev[7][97] & ~x[19];
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & x[28];
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & ~x[19];
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & ~x[49];
			partial_clause[8][12] 	= partial_clause_prev[8][12] & x[6];
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & ~x[48];
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & x[56];
			partial_clause[8][46] 	= partial_clause_prev[8][46] & ~x[45];
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & ~x[34];
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & ~x[29] & ~x[56];
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & ~x[28] & ~x[40] & ~x[56];
			partial_clause[8][57] 	= partial_clause_prev[8][57] & ~x[14];
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & ~x[57];
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & ~x[11] & ~x[41] & ~x[47];
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & ~x[57];
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & ~x[42];
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & ~x[28] & ~x[56];
			partial_clause[8][76] 	= partial_clause_prev[8][76] & ~x[18];
			partial_clause[8][77] 	= partial_clause_prev[8][77] & ~x[42];
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & ~x[29] & ~x[56];
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & ~x[29] & ~x[56];
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & ~x[29];
			partial_clause[8][89] 	= partial_clause_prev[8][89] & ~x[42] & ~x[57];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & ~x[46];
			partial_clause[8][92] 	= partial_clause_prev[8][92] & ~x[43];
			partial_clause[8][93] 	= partial_clause_prev[8][93] & ~x[46];
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & ~x[16] & ~x[28] & ~x[55];
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & x[33];
			partial_clause[9][4] 	= partial_clause_prev[9][4] & ~x[16];
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & ~x[1];
			partial_clause[9][11] 	= partial_clause_prev[9][11] & ~x[1];
			partial_clause[9][12] 	= partial_clause_prev[9][12] & ~x[13];
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & x[61];
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & 1'b1;
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & x[61];
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & x[53];
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & x[61];
			partial_clause[9][49] 	= partial_clause_prev[9][49] & x[61];
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & ~x[61] & ~x[62];
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & ~x[61];
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & ~x[26] & ~x[52];
			partial_clause[9][60] 	= partial_clause_prev[9][60] & ~x[14];
			partial_clause[9][61] 	= partial_clause_prev[9][61] & ~x[33];
			partial_clause[9][62] 	= partial_clause_prev[9][62] & ~x[16];
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & ~x[62];
			partial_clause[9][68] 	= partial_clause_prev[9][68] & ~x[21] & ~x[61];
			partial_clause[9][69] 	= partial_clause_prev[9][69] & ~x[17];
			partial_clause[9][70] 	= partial_clause_prev[9][70] & ~x[14];
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & ~x[14];
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & ~x[18];
			partial_clause[9][78] 	= partial_clause_prev[9][78] & ~x[26] & ~x[50] & ~x[51] & ~x[54];
			partial_clause[9][79] 	= partial_clause_prev[9][79] & ~x[61];
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & ~x[18] & ~x[43];
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & ~x[40];
			partial_clause[9][87] 	= partial_clause_prev[9][87] & ~x[24] & ~x[25] & ~x[26] & ~x[50];
			partial_clause[9][88] 	= partial_clause_prev[9][88] & ~x[52];
			partial_clause[9][89] 	= partial_clause_prev[9][89] & ~x[20];
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & ~x[46];
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & ~x[53] & ~x[54];
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
		end
	end
endmodule


module HCB_6 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & ~x[23] & ~x[50];
			partial_clause[0][1] 	= partial_clause_prev[0][1] & ~x[23];
			partial_clause[0][2] 	= partial_clause_prev[0][2] & ~x[51];
			partial_clause[0][3] 	= partial_clause_prev[0][3] & ~x[50];
			partial_clause[0][4] 	= partial_clause_prev[0][4] & ~x[21] & ~x[24];
			partial_clause[0][5] 	= partial_clause_prev[0][5] & ~x[21] & ~x[23] & ~x[24] & ~x[38];
			partial_clause[0][6] 	= partial_clause_prev[0][6] & ~x[23] & ~x[24];
			partial_clause[0][7] 	= partial_clause_prev[0][7] & ~x[22] & ~x[51];
			partial_clause[0][8] 	= partial_clause_prev[0][8] & ~x[22];
			partial_clause[0][9] 	= partial_clause_prev[0][9] & ~x[24] & ~x[51] & ~x[52];
			partial_clause[0][10] 	= partial_clause_prev[0][10] & ~x[23] & ~x[52];
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & ~x[22] & ~x[51];
			partial_clause[0][13] 	= partial_clause_prev[0][13] & ~x[21];
			partial_clause[0][14] 	= partial_clause_prev[0][14] & ~x[51];
			partial_clause[0][15] 	= partial_clause_prev[0][15] & ~x[22] & ~x[23] & ~x[50];
			partial_clause[0][16] 	= partial_clause_prev[0][16] & ~x[50];
			partial_clause[0][17] 	= partial_clause_prev[0][17] & ~x[50];
			partial_clause[0][18] 	= partial_clause_prev[0][18] & ~x[24] & ~x[50];
			partial_clause[0][19] 	= partial_clause_prev[0][19] & ~x[24] & ~x[48];
			partial_clause[0][20] 	= partial_clause_prev[0][20] & ~x[22] & ~x[49] & ~x[50];
			partial_clause[0][21] 	= partial_clause_prev[0][21] & ~x[22] & ~x[25];
			partial_clause[0][22] 	= partial_clause_prev[0][22] & ~x[49];
			partial_clause[0][23] 	= partial_clause_prev[0][23] & ~x[22] & ~x[24] & ~x[49];
			partial_clause[0][24] 	= partial_clause_prev[0][24] & ~x[24] & ~x[51];
			partial_clause[0][25] 	= partial_clause_prev[0][25] & ~x[21];
			partial_clause[0][26] 	= partial_clause_prev[0][26] & ~x[51] & ~x[52];
			partial_clause[0][27] 	= partial_clause_prev[0][27] & ~x[51] & ~x[52];
			partial_clause[0][28] 	= partial_clause_prev[0][28] & ~x[22];
			partial_clause[0][29] 	= partial_clause_prev[0][29] & ~x[50];
			partial_clause[0][30] 	= partial_clause_prev[0][30] & ~x[38];
			partial_clause[0][31] 	= partial_clause_prev[0][31] & ~x[22] & ~x[24] & ~x[50];
			partial_clause[0][32] 	= partial_clause_prev[0][32] & ~x[21] & ~x[49] & ~x[52];
			partial_clause[0][33] 	= partial_clause_prev[0][33] & ~x[23] & ~x[24] & ~x[51];
			partial_clause[0][34] 	= partial_clause_prev[0][34] & ~x[24];
			partial_clause[0][35] 	= partial_clause_prev[0][35] & ~x[24] & ~x[51] & ~x[52];
			partial_clause[0][36] 	= partial_clause_prev[0][36] & ~x[23] & ~x[50];
			partial_clause[0][37] 	= partial_clause_prev[0][37] & ~x[24] & ~x[25];
			partial_clause[0][38] 	= partial_clause_prev[0][38] & ~x[25];
			partial_clause[0][39] 	= partial_clause_prev[0][39] & ~x[52];
			partial_clause[0][40] 	= partial_clause_prev[0][40] & ~x[23] & ~x[50];
			partial_clause[0][41] 	= partial_clause_prev[0][41] & ~x[22] & ~x[24];
			partial_clause[0][42] 	= partial_clause_prev[0][42] & ~x[22] & ~x[52];
			partial_clause[0][43] 	= partial_clause_prev[0][43] & ~x[49] & ~x[51] & ~x[52];
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & ~x[24];
			partial_clause[0][46] 	= partial_clause_prev[0][46] & ~x[24] & ~x[52];
			partial_clause[0][47] 	= partial_clause_prev[0][47] & ~x[21] & ~x[24] & ~x[25];
			partial_clause[0][48] 	= partial_clause_prev[0][48] & ~x[24] & ~x[48] & ~x[52];
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & ~x[0] & ~x[2] & ~x[36];
			partial_clause[0][51] 	= partial_clause_prev[0][51] & ~x[1] & ~x[11] & x[51];
			partial_clause[0][52] 	= partial_clause_prev[0][52] & x[50];
			partial_clause[0][53] 	= partial_clause_prev[0][53] & ~x[6] & x[51];
			partial_clause[0][54] 	= partial_clause_prev[0][54] & ~x[31];
			partial_clause[0][55] 	= partial_clause_prev[0][55] & ~x[33] & x[50];
			partial_clause[0][56] 	= partial_clause_prev[0][56] & x[50];
			partial_clause[0][57] 	= partial_clause_prev[0][57] & x[22];
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & ~x[33] & ~x[40] & x[51];
			partial_clause[0][60] 	= partial_clause_prev[0][60] & x[50];
			partial_clause[0][61] 	= partial_clause_prev[0][61] & ~x[4] & ~x[37];
			partial_clause[0][62] 	= partial_clause_prev[0][62] & ~x[3] & ~x[4] & ~x[35] & x[51];
			partial_clause[0][63] 	= partial_clause_prev[0][63] & ~x[1] & ~x[32];
			partial_clause[0][64] 	= partial_clause_prev[0][64] & ~x[6];
			partial_clause[0][65] 	= partial_clause_prev[0][65] & x[51];
			partial_clause[0][66] 	= partial_clause_prev[0][66] & ~x[0] & ~x[3];
			partial_clause[0][67] 	= partial_clause_prev[0][67] & ~x[31];
			partial_clause[0][68] 	= partial_clause_prev[0][68] & x[23];
			partial_clause[0][69] 	= partial_clause_prev[0][69] & x[52];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & ~x[2] & ~x[4];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & ~x[3] & x[24];
			partial_clause[0][72] 	= partial_clause_prev[0][72] & x[51];
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & x[23];
			partial_clause[0][75] 	= partial_clause_prev[0][75] & ~x[11] & ~x[63];
			partial_clause[0][76] 	= partial_clause_prev[0][76] & ~x[3];
			partial_clause[0][77] 	= partial_clause_prev[0][77] & ~x[3] & ~x[7] & ~x[32];
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & ~x[0] & ~x[2] & ~x[9];
			partial_clause[0][81] 	= partial_clause_prev[0][81] & ~x[3];
			partial_clause[0][82] 	= partial_clause_prev[0][82] & ~x[39];
			partial_clause[0][83] 	= partial_clause_prev[0][83] & x[23] & ~x[38];
			partial_clause[0][84] 	= partial_clause_prev[0][84] & x[51];
			partial_clause[0][85] 	= partial_clause_prev[0][85] & ~x[10] & ~x[33];
			partial_clause[0][86] 	= partial_clause_prev[0][86] & ~x[3];
			partial_clause[0][87] 	= partial_clause_prev[0][87] & ~x[0] & ~x[31] & ~x[32];
			partial_clause[0][88] 	= partial_clause_prev[0][88] & ~x[2] & x[23];
			partial_clause[0][89] 	= partial_clause_prev[0][89] & ~x[0] & ~x[30];
			partial_clause[0][90] 	= partial_clause_prev[0][90] & ~x[0] & ~x[58];
			partial_clause[0][91] 	= partial_clause_prev[0][91] & x[23];
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & ~x[40] & x[51];
			partial_clause[0][94] 	= partial_clause_prev[0][94] & x[23];
			partial_clause[0][95] 	= partial_clause_prev[0][95] & ~x[3] & ~x[7];
			partial_clause[0][96] 	= partial_clause_prev[0][96] & ~x[0] & ~x[31];
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & ~x[14] & ~x[40];
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & ~x[28] & ~x[53];
			partial_clause[1][2] 	= partial_clause_prev[1][2] & ~x[27];
			partial_clause[1][3] 	= partial_clause_prev[1][3] & x[22] & ~x[55];
			partial_clause[1][4] 	= partial_clause_prev[1][4] & ~x[46];
			partial_clause[1][5] 	= partial_clause_prev[1][5] & x[22];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & ~x[10] & ~x[46] & ~x[53];
			partial_clause[1][7] 	= partial_clause_prev[1][7] & ~x[19] & ~x[55];
			partial_clause[1][8] 	= partial_clause_prev[1][8] & ~x[53];
			partial_clause[1][9] 	= partial_clause_prev[1][9] & x[22] & ~x[53];
			partial_clause[1][10] 	= partial_clause_prev[1][10] & ~x[18] & x[22];
			partial_clause[1][11] 	= partial_clause_prev[1][11] & ~x[26];
			partial_clause[1][12] 	= partial_clause_prev[1][12] & ~x[45] & ~x[53] & ~x[55];
			partial_clause[1][13] 	= partial_clause_prev[1][13] & ~x[18] & ~x[54];
			partial_clause[1][14] 	= partial_clause_prev[1][14] & x[22];
			partial_clause[1][15] 	= partial_clause_prev[1][15] & ~x[53];
			partial_clause[1][16] 	= partial_clause_prev[1][16] & ~x[26] & ~x[41];
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & ~x[0] & x[22];
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & x[50];
			partial_clause[1][23] 	= partial_clause_prev[1][23] & x[22] & ~x[53] & ~x[62];
			partial_clause[1][24] 	= partial_clause_prev[1][24] & ~x[18];
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & ~x[18] & x[50] & ~x[53];
			partial_clause[1][27] 	= partial_clause_prev[1][27] & x[22] & x[50] & ~x[53];
			partial_clause[1][28] 	= partial_clause_prev[1][28] & ~x[54];
			partial_clause[1][29] 	= partial_clause_prev[1][29] & x[50];
			partial_clause[1][30] 	= partial_clause_prev[1][30] & ~x[45];
			partial_clause[1][31] 	= partial_clause_prev[1][31] & ~x[18] & x[22];
			partial_clause[1][32] 	= partial_clause_prev[1][32] & ~x[53];
			partial_clause[1][33] 	= partial_clause_prev[1][33] & ~x[53];
			partial_clause[1][34] 	= partial_clause_prev[1][34] & ~x[55];
			partial_clause[1][35] 	= partial_clause_prev[1][35] & ~x[25] & x[50];
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & x[22] & ~x[53];
			partial_clause[1][38] 	= partial_clause_prev[1][38] & ~x[17] & x[22] & ~x[25];
			partial_clause[1][39] 	= partial_clause_prev[1][39] & x[22] & ~x[26] & x[50];
			partial_clause[1][40] 	= partial_clause_prev[1][40] & x[50] & ~x[53];
			partial_clause[1][41] 	= partial_clause_prev[1][41] & ~x[26] & ~x[27] & ~x[30];
			partial_clause[1][42] 	= partial_clause_prev[1][42] & ~x[25] & ~x[46];
			partial_clause[1][43] 	= partial_clause_prev[1][43] & ~x[17];
			partial_clause[1][44] 	= partial_clause_prev[1][44] & x[22] & ~x[26] & x[50];
			partial_clause[1][45] 	= partial_clause_prev[1][45] & ~x[19] & ~x[46] & x[50] & ~x[55];
			partial_clause[1][46] 	= partial_clause_prev[1][46] & x[22];
			partial_clause[1][47] 	= partial_clause_prev[1][47] & ~x[18] & ~x[25] & ~x[27] & ~x[45];
			partial_clause[1][48] 	= partial_clause_prev[1][48] & x[50] & ~x[54];
			partial_clause[1][49] 	= partial_clause_prev[1][49] & ~x[27];
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & ~x[37];
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & ~x[36] & x[54];
			partial_clause[1][56] 	= partial_clause_prev[1][56] & ~x[11];
			partial_clause[1][57] 	= partial_clause_prev[1][57] & ~x[37];
			partial_clause[1][58] 	= partial_clause_prev[1][58] & 1'b1;
			partial_clause[1][59] 	= partial_clause_prev[1][59] & x[26] & ~x[39];
			partial_clause[1][60] 	= partial_clause_prev[1][60] & ~x[7];
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & ~x[39];
			partial_clause[1][63] 	= partial_clause_prev[1][63] & ~x[11];
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & ~x[8] & ~x[37];
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & x[54] & ~x[63];
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & ~x[8] & ~x[38];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & x[25];
			partial_clause[1][77] 	= partial_clause_prev[1][77] & x[53];
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & ~x[35];
			partial_clause[1][81] 	= partial_clause_prev[1][81] & ~x[5];
			partial_clause[1][82] 	= partial_clause_prev[1][82] & ~x[35];
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & ~x[34];
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & ~x[9];
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & ~x[35];
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & ~x[12] & ~x[13];
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & ~x[14];
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & ~x[3] & ~x[30];
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & ~x[9];
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & ~x[31];
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & ~x[11] & ~x[33];
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & ~x[35];
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & ~x[60];
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & 1'b1;
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & ~x[11] & ~x[37] & ~x[60];
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & ~x[31];
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & ~x[4];
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & ~x[60];
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & ~x[60];
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & ~x[5];
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & ~x[38];
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & ~x[59];
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & ~x[5];
			partial_clause[2][96] 	= partial_clause_prev[2][96] & ~x[63];
			partial_clause[2][97] 	= partial_clause_prev[2][97] & ~x[10];
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & ~x[6];
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & ~x[43];
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & ~x[6];
			partial_clause[3][4] 	= partial_clause_prev[3][4] & ~x[3];
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & ~x[3];
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & ~x[3];
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & ~x[3];
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & ~x[13];
			partial_clause[3][18] 	= partial_clause_prev[3][18] & ~x[14];
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & ~x[8];
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & ~x[33];
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & ~x[39];
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & ~x[42];
			partial_clause[3][42] 	= partial_clause_prev[3][42] & ~x[7];
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & ~x[8];
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & ~x[14];
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & ~x[11];
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & ~x[36] & ~x[38];
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & ~x[63];
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & 1'b1;
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & ~x[10];
			partial_clause[3][68] 	= partial_clause_prev[3][68] & ~x[63];
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & ~x[36];
			partial_clause[3][77] 	= partial_clause_prev[3][77] & ~x[63];
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & ~x[62];
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & ~x[38];
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & ~x[40];
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & x[52];
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & x[17];
			partial_clause[4][8] 	= partial_clause_prev[4][8] & x[25] & x[52];
			partial_clause[4][9] 	= partial_clause_prev[4][9] & ~x[10];
			partial_clause[4][10] 	= partial_clause_prev[4][10] & ~x[37];
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & x[53];
			partial_clause[4][25] 	= partial_clause_prev[4][25] & x[53];
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & x[25];
			partial_clause[4][28] 	= partial_clause_prev[4][28] & x[53];
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & 1'b1;
			partial_clause[4][33] 	= partial_clause_prev[4][33] & x[25];
			partial_clause[4][34] 	= partial_clause_prev[4][34] & x[17];
			partial_clause[4][35] 	= partial_clause_prev[4][35] & x[53];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & x[52];
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & x[45];
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & ~x[10] & ~x[34];
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & ~x[3] & x[16];
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & 1'b1;
			partial_clause[4][50] 	= partial_clause_prev[4][50] & ~x[17] & ~x[45];
			partial_clause[4][51] 	= partial_clause_prev[4][51] & ~x[37];
			partial_clause[4][52] 	= partial_clause_prev[4][52] & ~x[12] & ~x[16] & ~x[17] & ~x[42] & ~x[43];
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & ~x[15] & ~x[17] & ~x[62];
			partial_clause[4][55] 	= partial_clause_prev[4][55] & ~x[60] & ~x[61];
			partial_clause[4][56] 	= partial_clause_prev[4][56] & ~x[43];
			partial_clause[4][57] 	= partial_clause_prev[4][57] & ~x[10] & ~x[15];
			partial_clause[4][58] 	= partial_clause_prev[4][58] & ~x[16] & ~x[17];
			partial_clause[4][59] 	= partial_clause_prev[4][59] & ~x[7] & ~x[35] & ~x[46];
			partial_clause[4][60] 	= partial_clause_prev[4][60] & ~x[6] & ~x[16] & ~x[18];
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & ~x[63];
			partial_clause[4][63] 	= partial_clause_prev[4][63] & ~x[17] & ~x[43];
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & ~x[8] & ~x[16];
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & ~x[46];
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & ~x[11] & ~x[45];
			partial_clause[4][72] 	= partial_clause_prev[4][72] & ~x[14] & ~x[16];
			partial_clause[4][73] 	= partial_clause_prev[4][73] & ~x[32] & ~x[37];
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & ~x[17] & ~x[42] & ~x[44];
			partial_clause[4][76] 	= partial_clause_prev[4][76] & ~x[4];
			partial_clause[4][77] 	= partial_clause_prev[4][77] & ~x[25] & ~x[35] & ~x[54];
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & ~x[14] & ~x[18];
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & ~x[16] & ~x[17] & ~x[18] & ~x[44];
			partial_clause[4][82] 	= partial_clause_prev[4][82] & ~x[44];
			partial_clause[4][83] 	= partial_clause_prev[4][83] & ~x[17] & ~x[42] & ~x[44];
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & ~x[16];
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & ~x[7];
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & ~x[5] & ~x[39];
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & ~x[39];
			partial_clause[4][94] 	= partial_clause_prev[4][94] & ~x[15];
			partial_clause[4][95] 	= partial_clause_prev[4][95] & ~x[45] & ~x[63];
			partial_clause[4][96] 	= partial_clause_prev[4][96] & ~x[37];
			partial_clause[4][97] 	= partial_clause_prev[4][97] & ~x[18] & ~x[44] & ~x[45] & ~x[63];
			partial_clause[4][98] 	= partial_clause_prev[4][98] & ~x[48];
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & ~x[0] & ~x[2] & ~x[30];
			partial_clause[5][1] 	= partial_clause_prev[5][1] & ~x[30];
			partial_clause[5][2] 	= partial_clause_prev[5][2] & ~x[2] & ~x[29];
			partial_clause[5][3] 	= partial_clause_prev[5][3] & ~x[39];
			partial_clause[5][4] 	= partial_clause_prev[5][4] & ~x[28];
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & ~x[30];
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & ~x[1];
			partial_clause[5][12] 	= partial_clause_prev[5][12] & ~x[2] & ~x[29];
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & ~x[4];
			partial_clause[5][19] 	= partial_clause_prev[5][19] & ~x[3];
			partial_clause[5][20] 	= partial_clause_prev[5][20] & ~x[1];
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & x[20];
			partial_clause[5][25] 	= partial_clause_prev[5][25] & ~x[1];
			partial_clause[5][26] 	= partial_clause_prev[5][26] & ~x[1];
			partial_clause[5][27] 	= partial_clause_prev[5][27] & ~x[7];
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & ~x[2];
			partial_clause[5][31] 	= partial_clause_prev[5][31] & ~x[2];
			partial_clause[5][32] 	= partial_clause_prev[5][32] & ~x[30];
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & ~x[2];
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & ~x[2] & ~x[3];
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & ~x[0] & ~x[56];
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & ~x[2];
			partial_clause[5][47] 	= partial_clause_prev[5][47] & ~x[58];
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & x[52];
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & x[24];
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & x[51];
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & x[51];
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & ~x[7];
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & ~x[11];
			partial_clause[5][91] 	= partial_clause_prev[5][91] & ~x[8] & x[24];
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & x[50];
			partial_clause[5][94] 	= partial_clause_prev[5][94] & ~x[37];
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & ~x[38];
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & ~x[8];
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & ~x[38];
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & ~x[40];
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & ~x[7];
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & ~x[37];
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & ~x[9];
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & ~x[9];
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & ~x[30];
			partial_clause[6][59] 	= partial_clause_prev[6][59] & ~x[7];
			partial_clause[6][60] 	= partial_clause_prev[6][60] & ~x[61];
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & ~x[46];
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & ~x[7];
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & ~x[3];
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & ~x[1] & ~x[3];
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & ~x[8];
			partial_clause[6][84] 	= partial_clause_prev[6][84] & ~x[4] & ~x[32];
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & ~x[31];
			partial_clause[6][89] 	= partial_clause_prev[6][89] & ~x[2] & ~x[3];
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & ~x[8];
			partial_clause[6][92] 	= partial_clause_prev[6][92] & ~x[5];
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & ~x[59];
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & ~x[32] & ~x[62];
			partial_clause[6][99] 	= partial_clause_prev[6][99] & ~x[4];
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & ~x[49];
			partial_clause[7][1] 	= partial_clause_prev[7][1] & ~x[19];
			partial_clause[7][2] 	= partial_clause_prev[7][2] & ~x[20];
			partial_clause[7][3] 	= partial_clause_prev[7][3] & ~x[47];
			partial_clause[7][4] 	= partial_clause_prev[7][4] & ~x[21];
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & ~x[21] & ~x[47];
			partial_clause[7][8] 	= partial_clause_prev[7][8] & ~x[48] & ~x[49];
			partial_clause[7][9] 	= partial_clause_prev[7][9] & ~x[20];
			partial_clause[7][10] 	= partial_clause_prev[7][10] & ~x[45];
			partial_clause[7][11] 	= partial_clause_prev[7][11] & ~x[47];
			partial_clause[7][12] 	= partial_clause_prev[7][12] & ~x[20];
			partial_clause[7][13] 	= partial_clause_prev[7][13] & ~x[21] & ~x[45] & ~x[46];
			partial_clause[7][14] 	= partial_clause_prev[7][14] & ~x[20] & ~x[46];
			partial_clause[7][15] 	= partial_clause_prev[7][15] & ~x[20] & ~x[21];
			partial_clause[7][16] 	= partial_clause_prev[7][16] & ~x[19] & ~x[21];
			partial_clause[7][17] 	= partial_clause_prev[7][17] & ~x[19] & ~x[21];
			partial_clause[7][18] 	= partial_clause_prev[7][18] & ~x[21] & ~x[46];
			partial_clause[7][19] 	= partial_clause_prev[7][19] & ~x[21];
			partial_clause[7][20] 	= partial_clause_prev[7][20] & ~x[49];
			partial_clause[7][21] 	= partial_clause_prev[7][21] & ~x[47] & ~x[48];
			partial_clause[7][22] 	= partial_clause_prev[7][22] & ~x[49];
			partial_clause[7][23] 	= partial_clause_prev[7][23] & ~x[37] & ~x[46];
			partial_clause[7][24] 	= partial_clause_prev[7][24] & ~x[19] & ~x[21] & ~x[47];
			partial_clause[7][25] 	= partial_clause_prev[7][25] & ~x[19] & ~x[21];
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & ~x[20] & ~x[42] & ~x[47];
			partial_clause[7][28] 	= partial_clause_prev[7][28] & ~x[49];
			partial_clause[7][29] 	= partial_clause_prev[7][29] & ~x[21] & ~x[47];
			partial_clause[7][30] 	= partial_clause_prev[7][30] & ~x[20] & ~x[47];
			partial_clause[7][31] 	= partial_clause_prev[7][31] & ~x[48];
			partial_clause[7][32] 	= partial_clause_prev[7][32] & ~x[21] & ~x[46];
			partial_clause[7][33] 	= partial_clause_prev[7][33] & ~x[20] & ~x[21] & ~x[48];
			partial_clause[7][34] 	= partial_clause_prev[7][34] & ~x[21] & ~x[47];
			partial_clause[7][35] 	= partial_clause_prev[7][35] & ~x[19] & ~x[47];
			partial_clause[7][36] 	= partial_clause_prev[7][36] & ~x[18] & ~x[21] & ~x[45];
			partial_clause[7][37] 	= partial_clause_prev[7][37] & ~x[21] & ~x[47];
			partial_clause[7][38] 	= partial_clause_prev[7][38] & ~x[47];
			partial_clause[7][39] 	= partial_clause_prev[7][39] & ~x[20] & ~x[46];
			partial_clause[7][40] 	= partial_clause_prev[7][40] & ~x[21] & ~x[45] & ~x[46];
			partial_clause[7][41] 	= partial_clause_prev[7][41] & ~x[48];
			partial_clause[7][42] 	= partial_clause_prev[7][42] & ~x[47];
			partial_clause[7][43] 	= partial_clause_prev[7][43] & ~x[5] & ~x[19] & ~x[44] & ~x[45];
			partial_clause[7][44] 	= partial_clause_prev[7][44] & ~x[21];
			partial_clause[7][45] 	= partial_clause_prev[7][45] & ~x[21] & ~x[47];
			partial_clause[7][46] 	= partial_clause_prev[7][46] & ~x[21] & ~x[47];
			partial_clause[7][47] 	= partial_clause_prev[7][47] & ~x[48];
			partial_clause[7][48] 	= partial_clause_prev[7][48] & ~x[45];
			partial_clause[7][49] 	= partial_clause_prev[7][49] & ~x[20] & ~x[48];
			partial_clause[7][50] 	= partial_clause_prev[7][50] & ~x[9];
			partial_clause[7][51] 	= partial_clause_prev[7][51] & ~x[37];
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & x[21];
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & ~x[38];
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & x[46];
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & ~x[11];
			partial_clause[7][82] 	= partial_clause_prev[7][82] & x[20];
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & ~x[12];
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & ~x[7];
			partial_clause[7][94] 	= partial_clause_prev[7][94] & x[20];
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & ~x[63];
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & x[49];
			partial_clause[8][1] 	= partial_clause_prev[8][1] & x[50];
			partial_clause[8][2] 	= partial_clause_prev[8][2] & ~x[12] & x[49];
			partial_clause[8][3] 	= partial_clause_prev[8][3] & ~x[44];
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & ~x[16] & x[21] & ~x[41];
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & ~x[43];
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & x[49];
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & ~x[43] & ~x[45];
			partial_clause[8][12] 	= partial_clause_prev[8][12] & ~x[14] & x[21] & ~x[43];
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & ~x[56];
			partial_clause[8][15] 	= partial_clause_prev[8][15] & ~x[40] & x[49];
			partial_clause[8][16] 	= partial_clause_prev[8][16] & ~x[40];
			partial_clause[8][17] 	= partial_clause_prev[8][17] & ~x[43] & ~x[44];
			partial_clause[8][18] 	= partial_clause_prev[8][18] & ~x[15] & ~x[17] & ~x[40] & ~x[43] & ~x[57];
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & ~x[14] & ~x[15] & ~x[34];
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & ~x[8] & ~x[10];
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & ~x[43];
			partial_clause[8][26] 	= partial_clause_prev[8][26] & x[23];
			partial_clause[8][27] 	= partial_clause_prev[8][27] & ~x[44];
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & x[23];
			partial_clause[8][30] 	= partial_clause_prev[8][30] & ~x[44];
			partial_clause[8][31] 	= partial_clause_prev[8][31] & x[49];
			partial_clause[8][32] 	= partial_clause_prev[8][32] & x[49];
			partial_clause[8][33] 	= partial_clause_prev[8][33] & ~x[43];
			partial_clause[8][34] 	= partial_clause_prev[8][34] & x[49];
			partial_clause[8][35] 	= partial_clause_prev[8][35] & ~x[31];
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & ~x[29] & ~x[58];
			partial_clause[8][38] 	= partial_clause_prev[8][38] & ~x[43] & ~x[44];
			partial_clause[8][39] 	= partial_clause_prev[8][39] & ~x[43];
			partial_clause[8][40] 	= partial_clause_prev[8][40] & x[23] & ~x[43];
			partial_clause[8][41] 	= partial_clause_prev[8][41] & x[22];
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & ~x[14] & ~x[34] & x[49];
			partial_clause[8][45] 	= partial_clause_prev[8][45] & ~x[43] & x[50] & ~x[56];
			partial_clause[8][46] 	= partial_clause_prev[8][46] & ~x[44] & x[49];
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & ~x[44];
			partial_clause[8][49] 	= partial_clause_prev[8][49] & ~x[15] & ~x[44] & x[49];
			partial_clause[8][50] 	= partial_clause_prev[8][50] & ~x[20] & ~x[48];
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & ~x[20] & ~x[22];
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & ~x[6];
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & ~x[21] & ~x[48];
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & ~x[20];
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & ~x[38] & ~x[39];
			partial_clause[8][63] 	= partial_clause_prev[8][63] & ~x[11];
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & ~x[20] & ~x[21];
			partial_clause[8][67] 	= partial_clause_prev[8][67] & ~x[20] & ~x[21];
			partial_clause[8][68] 	= partial_clause_prev[8][68] & ~x[10];
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & ~x[21] & ~x[48];
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & ~x[39] & ~x[48] & ~x[49];
			partial_clause[8][75] 	= partial_clause_prev[8][75] & ~x[8] & ~x[19] & ~x[62];
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & ~x[11];
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & ~x[9] & ~x[20] & ~x[35];
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & ~x[22];
			partial_clause[8][87] 	= partial_clause_prev[8][87] & ~x[20];
			partial_clause[8][88] 	= partial_clause_prev[8][88] & ~x[20];
			partial_clause[8][89] 	= partial_clause_prev[8][89] & ~x[20];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & ~x[20] & ~x[22];
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & ~x[48] & ~x[49];
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & ~x[19];
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & x[25];
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & x[25];
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & ~x[58];
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & x[25];
			partial_clause[9][7] 	= partial_clause_prev[9][7] & x[25];
			partial_clause[9][8] 	= partial_clause_prev[9][8] & x[25];
			partial_clause[9][9] 	= partial_clause_prev[9][9] & x[24];
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & x[25];
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & x[25];
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & x[46];
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & x[25];
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & x[25] & x[53];
			partial_clause[9][20] 	= partial_clause_prev[9][20] & x[25];
			partial_clause[9][21] 	= partial_clause_prev[9][21] & x[25] & ~x[58] & ~x[61];
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & x[25];
			partial_clause[9][26] 	= partial_clause_prev[9][26] & x[24];
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & x[25];
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & ~x[57];
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & x[25];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & x[25];
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & x[25];
			partial_clause[9][48] 	= partial_clause_prev[9][48] & ~x[60];
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & ~x[12];
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & ~x[39];
			partial_clause[9][59] 	= partial_clause_prev[9][59] & ~x[13];
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & ~x[12] & ~x[14] & ~x[16];
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & ~x[63];
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & ~x[40];
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & ~x[13] & ~x[15];
			partial_clause[9][88] 	= partial_clause_prev[9][88] & ~x[12] & ~x[15] & ~x[38];
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & ~x[15] & ~x[41] & ~x[62];
			partial_clause[9][99] 	= partial_clause_prev[9][99] & ~x[53];
		end
	end
endmodule


module HCB_7 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & ~x[14];
			partial_clause[0][1] 	= partial_clause_prev[0][1] & ~x[14] & ~x[41];
			partial_clause[0][2] 	= partial_clause_prev[0][2] & ~x[15] & ~x[41];
			partial_clause[0][3] 	= partial_clause_prev[0][3] & ~x[31] & ~x[40];
			partial_clause[0][4] 	= partial_clause_prev[0][4] & ~x[59];
			partial_clause[0][5] 	= partial_clause_prev[0][5] & ~x[40];
			partial_clause[0][6] 	= partial_clause_prev[0][6] & ~x[14] & ~x[30] & ~x[40];
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & ~x[14] & ~x[42];
			partial_clause[0][9] 	= partial_clause_prev[0][9] & ~x[14] & ~x[40];
			partial_clause[0][10] 	= partial_clause_prev[0][10] & ~x[14] & ~x[15];
			partial_clause[0][11] 	= partial_clause_prev[0][11] & ~x[14] & ~x[16];
			partial_clause[0][12] 	= partial_clause_prev[0][12] & ~x[16];
			partial_clause[0][13] 	= partial_clause_prev[0][13] & ~x[14] & ~x[15];
			partial_clause[0][14] 	= partial_clause_prev[0][14] & ~x[27] & ~x[31];
			partial_clause[0][15] 	= partial_clause_prev[0][15] & ~x[41];
			partial_clause[0][16] 	= partial_clause_prev[0][16] & ~x[14];
			partial_clause[0][17] 	= partial_clause_prev[0][17] & ~x[41];
			partial_clause[0][18] 	= partial_clause_prev[0][18] & ~x[15] & ~x[42];
			partial_clause[0][19] 	= partial_clause_prev[0][19] & ~x[13];
			partial_clause[0][20] 	= partial_clause_prev[0][20] & ~x[42];
			partial_clause[0][21] 	= partial_clause_prev[0][21] & ~x[42] & ~x[58];
			partial_clause[0][22] 	= partial_clause_prev[0][22] & ~x[41];
			partial_clause[0][23] 	= partial_clause_prev[0][23] & ~x[15] & ~x[41];
			partial_clause[0][24] 	= partial_clause_prev[0][24] & ~x[15];
			partial_clause[0][25] 	= partial_clause_prev[0][25] & ~x[13];
			partial_clause[0][26] 	= partial_clause_prev[0][26] & ~x[13];
			partial_clause[0][27] 	= partial_clause_prev[0][27] & ~x[15];
			partial_clause[0][28] 	= partial_clause_prev[0][28] & ~x[13] & ~x[42];
			partial_clause[0][29] 	= partial_clause_prev[0][29] & ~x[2] & ~x[16] & ~x[40];
			partial_clause[0][30] 	= partial_clause_prev[0][30] & ~x[13] & ~x[15];
			partial_clause[0][31] 	= partial_clause_prev[0][31] & ~x[13] & ~x[41];
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & ~x[13];
			partial_clause[0][34] 	= partial_clause_prev[0][34] & x[7];
			partial_clause[0][35] 	= partial_clause_prev[0][35] & ~x[41];
			partial_clause[0][36] 	= partial_clause_prev[0][36] & ~x[41] & ~x[59];
			partial_clause[0][37] 	= partial_clause_prev[0][37] & ~x[15] & ~x[41];
			partial_clause[0][38] 	= partial_clause_prev[0][38] & ~x[12] & ~x[14];
			partial_clause[0][39] 	= partial_clause_prev[0][39] & ~x[15] & ~x[41];
			partial_clause[0][40] 	= partial_clause_prev[0][40] & ~x[41] & ~x[43];
			partial_clause[0][41] 	= partial_clause_prev[0][41] & ~x[15] & ~x[54];
			partial_clause[0][42] 	= partial_clause_prev[0][42] & ~x[12];
			partial_clause[0][43] 	= partial_clause_prev[0][43] & ~x[12] & ~x[42];
			partial_clause[0][44] 	= partial_clause_prev[0][44] & ~x[16] & ~x[41];
			partial_clause[0][45] 	= partial_clause_prev[0][45] & ~x[13] & ~x[15] & ~x[42];
			partial_clause[0][46] 	= partial_clause_prev[0][46] & ~x[14] & ~x[16];
			partial_clause[0][47] 	= partial_clause_prev[0][47] & ~x[13];
			partial_clause[0][48] 	= partial_clause_prev[0][48] & ~x[14] & ~x[42];
			partial_clause[0][49] 	= partial_clause_prev[0][49] & ~x[14] & ~x[15] & ~x[41];
			partial_clause[0][50] 	= partial_clause_prev[0][50] & ~x[24];
			partial_clause[0][51] 	= partial_clause_prev[0][51] & ~x[1];
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & ~x[34] & ~x[62];
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & ~x[54] & ~x[58];
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & ~x[5] & ~x[24] & ~x[34] & ~x[36] & ~x[60];
			partial_clause[0][59] 	= partial_clause_prev[0][59] & ~x[30];
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & ~x[32] & ~x[35] & ~x[36];
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & ~x[58];
			partial_clause[0][65] 	= partial_clause_prev[0][65] & ~x[32];
			partial_clause[0][66] 	= partial_clause_prev[0][66] & ~x[58];
			partial_clause[0][67] 	= partial_clause_prev[0][67] & ~x[34] & ~x[36];
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & ~x[0] & ~x[55];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & ~x[0];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & ~x[4];
			partial_clause[0][73] 	= partial_clause_prev[0][73] & ~x[32] & ~x[62] & ~x[63];
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & ~x[33];
			partial_clause[0][76] 	= partial_clause_prev[0][76] & x[14];
			partial_clause[0][77] 	= partial_clause_prev[0][77] & ~x[26] & ~x[27];
			partial_clause[0][78] 	= partial_clause_prev[0][78] & ~x[56];
			partial_clause[0][79] 	= partial_clause_prev[0][79] & ~x[61] & ~x[63];
			partial_clause[0][80] 	= partial_clause_prev[0][80] & ~x[5] & ~x[33];
			partial_clause[0][81] 	= partial_clause_prev[0][81] & ~x[33] & ~x[63];
			partial_clause[0][82] 	= partial_clause_prev[0][82] & ~x[5] & ~x[35] & ~x[36] & ~x[37];
			partial_clause[0][83] 	= partial_clause_prev[0][83] & ~x[33];
			partial_clause[0][84] 	= partial_clause_prev[0][84] & ~x[2];
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & ~x[57] & ~x[61] & ~x[63];
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & ~x[2];
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & ~x[30];
			partial_clause[0][92] 	= partial_clause_prev[0][92] & ~x[31] & ~x[35];
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & 1'b1;
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & ~x[0] & ~x[1] & x[14];
			partial_clause[0][98] 	= partial_clause_prev[0][98] & ~x[8];
			partial_clause[0][99] 	= partial_clause_prev[0][99] & ~x[34] & ~x[62];
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[19];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & ~x[36];
			partial_clause[1][4] 	= partial_clause_prev[1][4] & ~x[47];
			partial_clause[1][5] 	= partial_clause_prev[1][5] & ~x[9] & ~x[17];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & ~x[3];
			partial_clause[1][9] 	= partial_clause_prev[1][9] & ~x[45];
			partial_clause[1][10] 	= partial_clause_prev[1][10] & ~x[17] & ~x[63];
			partial_clause[1][11] 	= partial_clause_prev[1][11] & ~x[46] & ~x[63];
			partial_clause[1][12] 	= partial_clause_prev[1][12] & ~x[63];
			partial_clause[1][13] 	= partial_clause_prev[1][13] & ~x[8];
			partial_clause[1][14] 	= partial_clause_prev[1][14] & ~x[45];
			partial_clause[1][15] 	= partial_clause_prev[1][15] & ~x[9] & ~x[45];
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & ~x[9] & ~x[45];
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & ~x[45] & ~x[47] & ~x[62];
			partial_clause[1][21] 	= partial_clause_prev[1][21] & ~x[17];
			partial_clause[1][22] 	= partial_clause_prev[1][22] & ~x[46];
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & ~x[8];
			partial_clause[1][25] 	= partial_clause_prev[1][25] & ~x[49];
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & ~x[32];
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & ~x[17];
			partial_clause[1][30] 	= partial_clause_prev[1][30] & ~x[17];
			partial_clause[1][31] 	= partial_clause_prev[1][31] & ~x[8];
			partial_clause[1][32] 	= partial_clause_prev[1][32] & ~x[17];
			partial_clause[1][33] 	= partial_clause_prev[1][33] & ~x[47];
			partial_clause[1][34] 	= partial_clause_prev[1][34] & ~x[45];
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & ~x[45];
			partial_clause[1][37] 	= partial_clause_prev[1][37] & ~x[45] & ~x[46] & ~x[63];
			partial_clause[1][38] 	= partial_clause_prev[1][38] & ~x[21] & ~x[46];
			partial_clause[1][39] 	= partial_clause_prev[1][39] & ~x[33] & ~x[46];
			partial_clause[1][40] 	= partial_clause_prev[1][40] & ~x[17] & ~x[63];
			partial_clause[1][41] 	= partial_clause_prev[1][41] & ~x[10];
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & ~x[36];
			partial_clause[1][45] 	= partial_clause_prev[1][45] & ~x[18];
			partial_clause[1][46] 	= partial_clause_prev[1][46] & ~x[17] & ~x[22];
			partial_clause[1][47] 	= partial_clause_prev[1][47] & ~x[9];
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & ~x[35] & ~x[63];
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & ~x[3];
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & ~x[27];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & ~x[30];
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & ~x[28];
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & x[18];
			partial_clause[1][74] 	= partial_clause_prev[1][74] & ~x[53];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & x[9];
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & ~x[41] & ~x[42];
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & x[46];
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & x[45];
			partial_clause[1][84] 	= partial_clause_prev[1][84] & x[48];
			partial_clause[1][85] 	= partial_clause_prev[1][85] & ~x[55];
			partial_clause[1][86] 	= partial_clause_prev[1][86] & ~x[29] & x[45];
			partial_clause[1][87] 	= partial_clause_prev[1][87] & ~x[0];
			partial_clause[1][88] 	= partial_clause_prev[1][88] & ~x[26];
			partial_clause[1][89] 	= partial_clause_prev[1][89] & ~x[42];
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & x[46];
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & ~x[14] & ~x[29];
			partial_clause[1][95] 	= partial_clause_prev[1][95] & ~x[0];
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & x[45];
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & ~x[26];
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & ~x[56];
			partial_clause[2][32] 	= partial_clause_prev[2][32] & ~x[27];
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & ~x[1];
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & ~x[55];
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & x[37];
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & ~x[23] & ~x[61];
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & ~x[63];
			partial_clause[2][53] 	= partial_clause_prev[2][53] & ~x[23] & ~x[51];
			partial_clause[2][54] 	= partial_clause_prev[2][54] & ~x[24] & ~x[51] & ~x[63];
			partial_clause[2][55] 	= partial_clause_prev[2][55] & ~x[30];
			partial_clause[2][56] 	= partial_clause_prev[2][56] & ~x[32];
			partial_clause[2][57] 	= partial_clause_prev[2][57] & ~x[24] & ~x[63];
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & ~x[62] & ~x[63];
			partial_clause[2][60] 	= partial_clause_prev[2][60] & ~x[25] & ~x[51] & ~x[62];
			partial_clause[2][61] 	= partial_clause_prev[2][61] & ~x[52] & ~x[62];
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & ~x[3] & ~x[4] & ~x[36];
			partial_clause[2][64] 	= partial_clause_prev[2][64] & ~x[26] & ~x[28];
			partial_clause[2][65] 	= partial_clause_prev[2][65] & ~x[51];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & ~x[51] & ~x[62];
			partial_clause[2][67] 	= partial_clause_prev[2][67] & ~x[3];
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & ~x[52];
			partial_clause[2][70] 	= partial_clause_prev[2][70] & ~x[63];
			partial_clause[2][71] 	= partial_clause_prev[2][71] & ~x[26] & ~x[27];
			partial_clause[2][72] 	= partial_clause_prev[2][72] & ~x[23] & ~x[59];
			partial_clause[2][73] 	= partial_clause_prev[2][73] & ~x[60];
			partial_clause[2][74] 	= partial_clause_prev[2][74] & ~x[35] & ~x[62] & ~x[63];
			partial_clause[2][75] 	= partial_clause_prev[2][75] & ~x[25] & ~x[26];
			partial_clause[2][76] 	= partial_clause_prev[2][76] & ~x[63];
			partial_clause[2][77] 	= partial_clause_prev[2][77] & ~x[53];
			partial_clause[2][78] 	= partial_clause_prev[2][78] & ~x[22];
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & ~x[24];
			partial_clause[2][81] 	= partial_clause_prev[2][81] & ~x[24] & ~x[50] & ~x[61];
			partial_clause[2][82] 	= partial_clause_prev[2][82] & ~x[53];
			partial_clause[2][83] 	= partial_clause_prev[2][83] & ~x[61];
			partial_clause[2][84] 	= partial_clause_prev[2][84] & ~x[36];
			partial_clause[2][85] 	= partial_clause_prev[2][85] & ~x[29] & ~x[62];
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & ~x[26] & ~x[52] & ~x[60];
			partial_clause[2][88] 	= partial_clause_prev[2][88] & ~x[24];
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & ~x[51];
			partial_clause[2][92] 	= partial_clause_prev[2][92] & ~x[53];
			partial_clause[2][93] 	= partial_clause_prev[2][93] & ~x[24] & ~x[61];
			partial_clause[2][94] 	= partial_clause_prev[2][94] & ~x[61];
			partial_clause[2][95] 	= partial_clause_prev[2][95] & ~x[50] & ~x[62];
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & ~x[63];
			partial_clause[2][98] 	= partial_clause_prev[2][98] & ~x[25];
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & ~x[37] & ~x[39];
			partial_clause[3][1] 	= partial_clause_prev[3][1] & ~x[41];
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & ~x[39] & ~x[41] & ~x[42];
			partial_clause[3][4] 	= partial_clause_prev[3][4] & ~x[38] & ~x[40];
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & ~x[38] & ~x[41];
			partial_clause[3][7] 	= partial_clause_prev[3][7] & ~x[38] & ~x[41];
			partial_clause[3][8] 	= partial_clause_prev[3][8] & ~x[25];
			partial_clause[3][9] 	= partial_clause_prev[3][9] & ~x[38];
			partial_clause[3][10] 	= partial_clause_prev[3][10] & ~x[36] & ~x[39];
			partial_clause[3][11] 	= partial_clause_prev[3][11] & ~x[36];
			partial_clause[3][12] 	= partial_clause_prev[3][12] & ~x[36];
			partial_clause[3][13] 	= partial_clause_prev[3][13] & ~x[24];
			partial_clause[3][14] 	= partial_clause_prev[3][14] & ~x[38];
			partial_clause[3][15] 	= partial_clause_prev[3][15] & ~x[37] & ~x[39];
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & ~x[36] & ~x[42];
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & ~x[3] & ~x[38] & ~x[41];
			partial_clause[3][21] 	= partial_clause_prev[3][21] & ~x[2] & ~x[37] & ~x[39];
			partial_clause[3][22] 	= partial_clause_prev[3][22] & ~x[39] & ~x[41];
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & ~x[41] & ~x[42];
			partial_clause[3][25] 	= partial_clause_prev[3][25] & ~x[41];
			partial_clause[3][26] 	= partial_clause_prev[3][26] & ~x[40] & ~x[41] & ~x[42];
			partial_clause[3][27] 	= partial_clause_prev[3][27] & ~x[37] & ~x[42];
			partial_clause[3][28] 	= partial_clause_prev[3][28] & ~x[0] & ~x[6] & ~x[38];
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & ~x[36] & ~x[39] & ~x[40];
			partial_clause[3][31] 	= partial_clause_prev[3][31] & ~x[40];
			partial_clause[3][32] 	= partial_clause_prev[3][32] & ~x[38];
			partial_clause[3][33] 	= partial_clause_prev[3][33] & ~x[38];
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & ~x[38];
			partial_clause[3][37] 	= partial_clause_prev[3][37] & ~x[38];
			partial_clause[3][38] 	= partial_clause_prev[3][38] & ~x[1] & ~x[38];
			partial_clause[3][39] 	= partial_clause_prev[3][39] & ~x[38];
			partial_clause[3][40] 	= partial_clause_prev[3][40] & ~x[37] & ~x[39];
			partial_clause[3][41] 	= partial_clause_prev[3][41] & ~x[37];
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & ~x[7] & ~x[39] & ~x[42];
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & ~x[41];
			partial_clause[3][46] 	= partial_clause_prev[3][46] & ~x[39] & ~x[41];
			partial_clause[3][47] 	= partial_clause_prev[3][47] & ~x[37] & ~x[39] & ~x[42];
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & ~x[38] & ~x[41] & ~x[42];
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & ~x[1] & x[42];
			partial_clause[3][53] 	= partial_clause_prev[3][53] & ~x[54];
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & x[40];
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & ~x[30];
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & ~x[26] & x[40];
			partial_clause[3][62] 	= partial_clause_prev[3][62] & ~x[58];
			partial_clause[3][63] 	= partial_clause_prev[3][63] & ~x[31];
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & 1'b1;
			partial_clause[3][66] 	= partial_clause_prev[3][66] & ~x[25];
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & ~x[30];
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & x[42];
			partial_clause[3][74] 	= partial_clause_prev[3][74] & x[14];
			partial_clause[3][75] 	= partial_clause_prev[3][75] & ~x[31];
			partial_clause[3][76] 	= partial_clause_prev[3][76] & ~x[3];
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & ~x[59];
			partial_clause[3][81] 	= partial_clause_prev[3][81] & x[41];
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & ~x[31];
			partial_clause[3][85] 	= partial_clause_prev[3][85] & ~x[28] & ~x[59];
			partial_clause[3][86] 	= partial_clause_prev[3][86] & ~x[31];
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & x[14];
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & ~x[4];
			partial_clause[3][94] 	= partial_clause_prev[3][94] & ~x[58];
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & ~x[60];
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & x[15];
			partial_clause[4][7] 	= partial_clause_prev[4][7] & x[16];
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & x[16];
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & x[16];
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & ~x[26];
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & x[16];
			partial_clause[4][20] 	= partial_clause_prev[4][20] & ~x[51];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & ~x[24];
			partial_clause[4][22] 	= partial_clause_prev[4][22] & x[16] & ~x[54];
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & ~x[26];
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & 1'b1;
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & ~x[2];
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & x[15];
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & 1'b1;
			partial_clause[4][50] 	= partial_clause_prev[4][50] & ~x[8];
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & ~x[7];
			partial_clause[4][58] 	= partial_clause_prev[4][58] & ~x[0];
			partial_clause[4][59] 	= partial_clause_prev[4][59] & ~x[1] & ~x[10];
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & ~x[52];
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & ~x[29];
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & ~x[28];
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & ~x[58];
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & ~x[30];
			partial_clause[4][74] 	= partial_clause_prev[4][74] & ~x[3];
			partial_clause[4][75] 	= partial_clause_prev[4][75] & ~x[31];
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & ~x[15];
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & ~x[25];
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & ~x[28];
			partial_clause[4][83] 	= partial_clause_prev[4][83] & ~x[28];
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & ~x[28];
			partial_clause[4][87] 	= partial_clause_prev[4][87] & ~x[55];
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & ~x[29];
			partial_clause[4][92] 	= partial_clause_prev[4][92] & ~x[8];
			partial_clause[4][93] 	= partial_clause_prev[4][93] & ~x[16];
			partial_clause[4][94] 	= partial_clause_prev[4][94] & ~x[57];
			partial_clause[4][95] 	= partial_clause_prev[4][95] & ~x[8];
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & ~x[0] & ~x[39];
			partial_clause[4][99] 	= partial_clause_prev[4][99] & ~x[0];
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & ~x[22];
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & ~x[23];
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & ~x[39];
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & ~x[39];
			partial_clause[5][17] 	= partial_clause_prev[5][17] & ~x[38] & ~x[41];
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & ~x[29];
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & ~x[39];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & ~x[39];
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & ~x[37] & ~x[39];
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & ~x[39];
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & ~x[41];
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & ~x[38];
			partial_clause[5][36] 	= partial_clause_prev[5][36] & ~x[41];
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & ~x[41];
			partial_clause[5][41] 	= partial_clause_prev[5][41] & ~x[38];
			partial_clause[5][42] 	= partial_clause_prev[5][42] & ~x[41];
			partial_clause[5][43] 	= partial_clause_prev[5][43] & ~x[26];
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & ~x[38];
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & x[42];
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & ~x[3];
			partial_clause[5][54] 	= partial_clause_prev[5][54] & x[13];
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & ~x[56];
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & x[14];
			partial_clause[5][61] 	= partial_clause_prev[5][61] & ~x[61];
			partial_clause[5][62] 	= partial_clause_prev[5][62] & x[14];
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & ~x[54];
			partial_clause[5][65] 	= partial_clause_prev[5][65] & ~x[2];
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & x[14];
			partial_clause[5][69] 	= partial_clause_prev[5][69] & ~x[55];
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & ~x[28];
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & ~x[26];
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & x[41];
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & ~x[58];
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & x[14];
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & ~x[0] & ~x[56];
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & ~x[1];
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & ~x[28];
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & ~x[58];
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & ~x[61];
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & ~x[32];
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & ~x[30] & x[38];
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & ~x[59];
			partial_clause[6][39] 	= partial_clause_prev[6][39] & ~x[0];
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & ~x[32];
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & ~x[30];
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & ~x[38];
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & ~x[23];
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & ~x[1];
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & ~x[38];
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & ~x[38];
			partial_clause[6][75] 	= partial_clause_prev[6][75] & ~x[54];
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & ~x[53];
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & ~x[37];
			partial_clause[6][82] 	= partial_clause_prev[6][82] & ~x[25] & ~x[59];
			partial_clause[6][83] 	= partial_clause_prev[6][83] & ~x[30];
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & ~x[38];
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & ~x[59];
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & ~x[37];
			partial_clause[6][96] 	= partial_clause_prev[6][96] & ~x[59];
			partial_clause[6][97] 	= partial_clause_prev[6][97] & ~x[2];
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & ~x[23];
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & ~x[12] & ~x[63];
			partial_clause[7][1] 	= partial_clause_prev[7][1] & ~x[9] & ~x[10] & ~x[11] & ~x[63];
			partial_clause[7][2] 	= partial_clause_prev[7][2] & ~x[38] & ~x[62];
			partial_clause[7][3] 	= partial_clause_prev[7][3] & ~x[9];
			partial_clause[7][4] 	= partial_clause_prev[7][4] & ~x[10] & ~x[12] & ~x[38];
			partial_clause[7][5] 	= partial_clause_prev[7][5] & ~x[8] & ~x[61] & ~x[63];
			partial_clause[7][6] 	= partial_clause_prev[7][6] & ~x[11];
			partial_clause[7][7] 	= partial_clause_prev[7][7] & ~x[39] & ~x[62];
			partial_clause[7][8] 	= partial_clause_prev[7][8] & ~x[12] & ~x[49];
			partial_clause[7][9] 	= partial_clause_prev[7][9] & ~x[11] & ~x[12];
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & ~x[38];
			partial_clause[7][12] 	= partial_clause_prev[7][12] & ~x[10] & ~x[36] & ~x[51];
			partial_clause[7][13] 	= partial_clause_prev[7][13] & ~x[30] & ~x[62];
			partial_clause[7][14] 	= partial_clause_prev[7][14] & ~x[10] & ~x[49];
			partial_clause[7][15] 	= partial_clause_prev[7][15] & ~x[9];
			partial_clause[7][16] 	= partial_clause_prev[7][16] & ~x[11];
			partial_clause[7][17] 	= partial_clause_prev[7][17] & ~x[38];
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & ~x[11];
			partial_clause[7][20] 	= partial_clause_prev[7][20] & ~x[37] & ~x[38];
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & ~x[11];
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & ~x[38];
			partial_clause[7][25] 	= partial_clause_prev[7][25] & ~x[34] & ~x[51];
			partial_clause[7][26] 	= partial_clause_prev[7][26] & ~x[12];
			partial_clause[7][27] 	= partial_clause_prev[7][27] & ~x[8];
			partial_clause[7][28] 	= partial_clause_prev[7][28] & ~x[12] & ~x[32];
			partial_clause[7][29] 	= partial_clause_prev[7][29] & ~x[11] & ~x[36] & ~x[38];
			partial_clause[7][30] 	= partial_clause_prev[7][30] & ~x[10] & ~x[51];
			partial_clause[7][31] 	= partial_clause_prev[7][31] & ~x[4] & ~x[11] & ~x[61];
			partial_clause[7][32] 	= partial_clause_prev[7][32] & ~x[35];
			partial_clause[7][33] 	= partial_clause_prev[7][33] & ~x[10];
			partial_clause[7][34] 	= partial_clause_prev[7][34] & ~x[10];
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & ~x[35];
			partial_clause[7][37] 	= partial_clause_prev[7][37] & ~x[38];
			partial_clause[7][38] 	= partial_clause_prev[7][38] & ~x[10] & ~x[38];
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & ~x[37];
			partial_clause[7][42] 	= partial_clause_prev[7][42] & ~x[36] & ~x[39];
			partial_clause[7][43] 	= partial_clause_prev[7][43] & ~x[34];
			partial_clause[7][44] 	= partial_clause_prev[7][44] & ~x[12] & ~x[34] & ~x[61];
			partial_clause[7][45] 	= partial_clause_prev[7][45] & ~x[8];
			partial_clause[7][46] 	= partial_clause_prev[7][46] & ~x[12] & ~x[36] & ~x[62];
			partial_clause[7][47] 	= partial_clause_prev[7][47] & ~x[10] & ~x[38];
			partial_clause[7][48] 	= partial_clause_prev[7][48] & ~x[7];
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & ~x[26];
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & ~x[1];
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & ~x[28];
			partial_clause[7][78] 	= partial_clause_prev[7][78] & ~x[29];
			partial_clause[7][79] 	= partial_clause_prev[7][79] & ~x[0];
			partial_clause[7][80] 	= partial_clause_prev[7][80] & ~x[53];
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & ~x[55] & ~x[61];
			partial_clause[8][1] 	= partial_clause_prev[8][1] & ~x[0] & ~x[6];
			partial_clause[8][2] 	= partial_clause_prev[8][2] & ~x[20] & x[40] & ~x[57];
			partial_clause[8][3] 	= partial_clause_prev[8][3] & ~x[3] & ~x[6] & x[12] & x[39];
			partial_clause[8][4] 	= partial_clause_prev[8][4] & ~x[6] & ~x[7] & x[40];
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & ~x[7] & x[39];
			partial_clause[8][9] 	= partial_clause_prev[8][9] & ~x[29];
			partial_clause[8][10] 	= partial_clause_prev[8][10] & ~x[29];
			partial_clause[8][11] 	= partial_clause_prev[8][11] & x[12] & ~x[62];
			partial_clause[8][12] 	= partial_clause_prev[8][12] & ~x[4];
			partial_clause[8][13] 	= partial_clause_prev[8][13] & ~x[7];
			partial_clause[8][14] 	= partial_clause_prev[8][14] & x[13];
			partial_clause[8][15] 	= partial_clause_prev[8][15] & x[39];
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & x[12] & ~x[27];
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & ~x[3];
			partial_clause[8][20] 	= partial_clause_prev[8][20] & ~x[4] & ~x[8] & x[40];
			partial_clause[8][21] 	= partial_clause_prev[8][21] & ~x[33];
			partial_clause[8][22] 	= partial_clause_prev[8][22] & ~x[7];
			partial_clause[8][23] 	= partial_clause_prev[8][23] & ~x[6] & ~x[26] & x[39];
			partial_clause[8][24] 	= partial_clause_prev[8][24] & x[39];
			partial_clause[8][25] 	= partial_clause_prev[8][25] & x[39];
			partial_clause[8][26] 	= partial_clause_prev[8][26] & x[40];
			partial_clause[8][27] 	= partial_clause_prev[8][27] & x[39] & ~x[50];
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & ~x[25];
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & ~x[61];
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & ~x[5] & ~x[7] & ~x[59];
			partial_clause[8][37] 	= partial_clause_prev[8][37] & ~x[6];
			partial_clause[8][38] 	= partial_clause_prev[8][38] & x[40] & ~x[56];
			partial_clause[8][39] 	= partial_clause_prev[8][39] & x[40];
			partial_clause[8][40] 	= partial_clause_prev[8][40] & ~x[52];
			partial_clause[8][41] 	= partial_clause_prev[8][41] & x[39];
			partial_clause[8][42] 	= partial_clause_prev[8][42] & ~x[2] & ~x[58];
			partial_clause[8][43] 	= partial_clause_prev[8][43] & ~x[6];
			partial_clause[8][44] 	= partial_clause_prev[8][44] & x[39];
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & x[39];
			partial_clause[8][49] 	= partial_clause_prev[8][49] & x[39];
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & ~x[11] & ~x[13] & ~x[27];
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & ~x[39] & ~x[40];
			partial_clause[8][59] 	= partial_clause_prev[8][59] & ~x[54];
			partial_clause[8][60] 	= partial_clause_prev[8][60] & ~x[10] & ~x[13];
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & ~x[28] & ~x[58];
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & ~x[37] & ~x[40] & ~x[59];
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & ~x[11] & ~x[12] & ~x[13] & ~x[30];
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & ~x[3];
			partial_clause[8][76] 	= partial_clause_prev[8][76] & ~x[30];
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & ~x[1];
			partial_clause[8][79] 	= partial_clause_prev[8][79] & ~x[31] & ~x[55];
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & ~x[3];
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & ~x[3];
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & ~x[0];
			partial_clause[8][96] 	= partial_clause_prev[8][96] & ~x[3] & ~x[38] & ~x[39] & ~x[40];
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & ~x[27];
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & ~x[21] & ~x[48];
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & ~x[50];
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & ~x[49];
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & ~x[3];
			partial_clause[9][12] 	= partial_clause_prev[9][12] & x[16] & ~x[50];
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & ~x[20];
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & ~x[23] & ~x[30];
			partial_clause[9][29] 	= partial_clause_prev[9][29] & ~x[20];
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & ~x[48];
			partial_clause[9][33] 	= partial_clause_prev[9][33] & ~x[21];
			partial_clause[9][34] 	= partial_clause_prev[9][34] & ~x[51];
			partial_clause[9][35] 	= partial_clause_prev[9][35] & 1'b1;
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & ~x[61];
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & ~x[51];
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & ~x[49];
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & ~x[3];
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & ~x[0];
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & ~x[57];
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
		end
	end
endmodule


module HCB_8 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & ~x[18];
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & x[56];
			partial_clause[0][4] 	= partial_clause_prev[0][4] & ~x[23];
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & x[0];
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & x[27];
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & ~x[21];
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & ~x[17];
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & ~x[19];
			partial_clause[0][34] 	= partial_clause_prev[0][34] & ~x[18];
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & ~x[51];
			partial_clause[0][52] 	= partial_clause_prev[0][52] & ~x[22];
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & ~x[28] & ~x[29];
			partial_clause[0][55] 	= partial_clause_prev[0][55] & ~x[18];
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & ~x[22];
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & ~x[1];
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & ~x[0] & ~x[16];
			partial_clause[0][76] 	= partial_clause_prev[0][76] & ~x[22];
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & ~x[29] & ~x[55];
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & ~x[0] & ~x[47];
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & ~x[22];
			partial_clause[0][86] 	= partial_clause_prev[0][86] & ~x[29];
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & ~x[1];
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & ~x[18];
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & ~x[50];
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & ~x[28] & ~x[29];
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & ~x[9] & ~x[38] & ~x[40];
			partial_clause[1][2] 	= partial_clause_prev[1][2] & ~x[9];
			partial_clause[1][3] 	= partial_clause_prev[1][3] & ~x[27] & ~x[39];
			partial_clause[1][4] 	= partial_clause_prev[1][4] & ~x[11] & ~x[54];
			partial_clause[1][5] 	= partial_clause_prev[1][5] & ~x[38];
			partial_clause[1][6] 	= partial_clause_prev[1][6] & ~x[9];
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & ~x[9];
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & ~x[10];
			partial_clause[1][12] 	= partial_clause_prev[1][12] & ~x[14] & ~x[28];
			partial_clause[1][13] 	= partial_clause_prev[1][13] & ~x[12] & ~x[38];
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & ~x[43];
			partial_clause[1][17] 	= partial_clause_prev[1][17] & ~x[38];
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & ~x[10];
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & ~x[0];
			partial_clause[1][28] 	= partial_clause_prev[1][28] & ~x[10];
			partial_clause[1][29] 	= partial_clause_prev[1][29] & ~x[27] & ~x[38];
			partial_clause[1][30] 	= partial_clause_prev[1][30] & ~x[10];
			partial_clause[1][31] 	= partial_clause_prev[1][31] & ~x[37];
			partial_clause[1][32] 	= partial_clause_prev[1][32] & ~x[27] & ~x[38];
			partial_clause[1][33] 	= partial_clause_prev[1][33] & ~x[27];
			partial_clause[1][34] 	= partial_clause_prev[1][34] & ~x[38];
			partial_clause[1][35] 	= partial_clause_prev[1][35] & ~x[10];
			partial_clause[1][36] 	= partial_clause_prev[1][36] & ~x[39];
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & ~x[10];
			partial_clause[1][43] 	= partial_clause_prev[1][43] & ~x[27];
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & ~x[42];
			partial_clause[1][47] 	= partial_clause_prev[1][47] & ~x[10];
			partial_clause[1][48] 	= partial_clause_prev[1][48] & ~x[0] & ~x[25];
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & x[37];
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & x[39] & ~x[50];
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & x[38];
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & ~x[46] & ~x[49];
			partial_clause[1][58] 	= partial_clause_prev[1][58] & ~x[21];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & x[38];
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & x[38];
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & ~x[50];
			partial_clause[1][74] 	= partial_clause_prev[1][74] & ~x[48];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & ~x[20];
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & ~x[48];
			partial_clause[1][82] 	= partial_clause_prev[1][82] & ~x[22] & ~x[48];
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & x[37];
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & ~x[4];
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & ~x[47];
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & ~x[19] & ~x[48];
			partial_clause[1][97] 	= partial_clause_prev[1][97] & ~x[47];
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & x[56];
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & x[58];
			partial_clause[2][7] 	= partial_clause_prev[2][7] & x[58];
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & x[56];
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & x[29];
			partial_clause[2][14] 	= partial_clause_prev[2][14] & x[1];
			partial_clause[2][15] 	= partial_clause_prev[2][15] & x[56];
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & x[56];
			partial_clause[2][19] 	= partial_clause_prev[2][19] & ~x[50];
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & x[58];
			partial_clause[2][22] 	= partial_clause_prev[2][22] & x[58];
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & x[40];
			partial_clause[2][25] 	= partial_clause_prev[2][25] & x[56];
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & x[57];
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & x[7];
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & ~x[2];
			partial_clause[2][51] 	= partial_clause_prev[2][51] & ~x[13] & ~x[40];
			partial_clause[2][52] 	= partial_clause_prev[2][52] & ~x[28];
			partial_clause[2][53] 	= partial_clause_prev[2][53] & ~x[14] & ~x[28] & ~x[41] & ~x[56];
			partial_clause[2][54] 	= partial_clause_prev[2][54] & ~x[41];
			partial_clause[2][55] 	= partial_clause_prev[2][55] & ~x[4] & ~x[16];
			partial_clause[2][56] 	= partial_clause_prev[2][56] & ~x[15];
			partial_clause[2][57] 	= partial_clause_prev[2][57] & ~x[14] & ~x[54];
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & ~x[13];
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & ~x[14] & ~x[26] & ~x[27];
			partial_clause[2][62] 	= partial_clause_prev[2][62] & ~x[15] & ~x[25] & ~x[29];
			partial_clause[2][63] 	= partial_clause_prev[2][63] & ~x[15];
			partial_clause[2][64] 	= partial_clause_prev[2][64] & ~x[43];
			partial_clause[2][65] 	= partial_clause_prev[2][65] & ~x[30];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & ~x[42] & ~x[55];
			partial_clause[2][67] 	= partial_clause_prev[2][67] & ~x[16];
			partial_clause[2][68] 	= partial_clause_prev[2][68] & ~x[15];
			partial_clause[2][69] 	= partial_clause_prev[2][69] & ~x[52];
			partial_clause[2][70] 	= partial_clause_prev[2][70] & ~x[14] & ~x[16];
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & ~x[14] & ~x[27];
			partial_clause[2][73] 	= partial_clause_prev[2][73] & ~x[13] & ~x[26] & ~x[29];
			partial_clause[2][74] 	= partial_clause_prev[2][74] & ~x[30] & ~x[43] & ~x[47];
			partial_clause[2][75] 	= partial_clause_prev[2][75] & ~x[2];
			partial_clause[2][76] 	= partial_clause_prev[2][76] & ~x[42] & ~x[57];
			partial_clause[2][77] 	= partial_clause_prev[2][77] & ~x[4];
			partial_clause[2][78] 	= partial_clause_prev[2][78] & ~x[15] & ~x[25] & ~x[50];
			partial_clause[2][79] 	= partial_clause_prev[2][79] & ~x[15] & ~x[44];
			partial_clause[2][80] 	= partial_clause_prev[2][80] & ~x[16] & ~x[43] & ~x[57];
			partial_clause[2][81] 	= partial_clause_prev[2][81] & ~x[1] & ~x[14] & ~x[41];
			partial_clause[2][82] 	= partial_clause_prev[2][82] & ~x[27] & ~x[40] & ~x[41];
			partial_clause[2][83] 	= partial_clause_prev[2][83] & ~x[14] & ~x[55];
			partial_clause[2][84] 	= partial_clause_prev[2][84] & ~x[15] & ~x[41];
			partial_clause[2][85] 	= partial_clause_prev[2][85] & ~x[15];
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & ~x[27] & ~x[54];
			partial_clause[2][88] 	= partial_clause_prev[2][88] & ~x[15];
			partial_clause[2][89] 	= partial_clause_prev[2][89] & ~x[24];
			partial_clause[2][90] 	= partial_clause_prev[2][90] & ~x[31] & ~x[42] & ~x[45];
			partial_clause[2][91] 	= partial_clause_prev[2][91] & ~x[26] & ~x[27] & ~x[57];
			partial_clause[2][92] 	= partial_clause_prev[2][92] & ~x[29] & ~x[53];
			partial_clause[2][93] 	= partial_clause_prev[2][93] & ~x[25] & ~x[42] & ~x[58];
			partial_clause[2][94] 	= partial_clause_prev[2][94] & ~x[16] & ~x[27];
			partial_clause[2][95] 	= partial_clause_prev[2][95] & ~x[13] & ~x[15] & ~x[16];
			partial_clause[2][96] 	= partial_clause_prev[2][96] & ~x[16] & ~x[23];
			partial_clause[2][97] 	= partial_clause_prev[2][97] & ~x[16] & ~x[29];
			partial_clause[2][98] 	= partial_clause_prev[2][98] & ~x[45];
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & ~x[4] & ~x[6];
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & ~x[4] & ~x[5] & ~x[17];
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & ~x[5];
			partial_clause[3][5] 	= partial_clause_prev[3][5] & ~x[2] & ~x[4] & ~x[5] & ~x[6];
			partial_clause[3][6] 	= partial_clause_prev[3][6] & ~x[7];
			partial_clause[3][7] 	= partial_clause_prev[3][7] & ~x[3];
			partial_clause[3][8] 	= partial_clause_prev[3][8] & ~x[5];
			partial_clause[3][9] 	= partial_clause_prev[3][9] & ~x[5] & ~x[6];
			partial_clause[3][10] 	= partial_clause_prev[3][10] & ~x[6] & ~x[47];
			partial_clause[3][11] 	= partial_clause_prev[3][11] & ~x[1] & ~x[3] & ~x[6];
			partial_clause[3][12] 	= partial_clause_prev[3][12] & ~x[3] & ~x[6];
			partial_clause[3][13] 	= partial_clause_prev[3][13] & ~x[2] & ~x[4] & ~x[6];
			partial_clause[3][14] 	= partial_clause_prev[3][14] & ~x[2] & ~x[4] & ~x[5];
			partial_clause[3][15] 	= partial_clause_prev[3][15] & ~x[5] & ~x[6];
			partial_clause[3][16] 	= partial_clause_prev[3][16] & ~x[3] & ~x[4] & ~x[5];
			partial_clause[3][17] 	= partial_clause_prev[3][17] & ~x[3] & ~x[4] & ~x[33] & ~x[46];
			partial_clause[3][18] 	= partial_clause_prev[3][18] & ~x[2] & ~x[6];
			partial_clause[3][19] 	= partial_clause_prev[3][19] & ~x[3];
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & ~x[4] & ~x[6] & ~x[21];
			partial_clause[3][22] 	= partial_clause_prev[3][22] & ~x[5];
			partial_clause[3][23] 	= partial_clause_prev[3][23] & ~x[2] & ~x[5] & ~x[49];
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & ~x[1];
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & ~x[3];
			partial_clause[3][28] 	= partial_clause_prev[3][28] & ~x[5];
			partial_clause[3][29] 	= partial_clause_prev[3][29] & ~x[3] & ~x[6];
			partial_clause[3][30] 	= partial_clause_prev[3][30] & ~x[2] & ~x[6];
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & ~x[2] & ~x[5] & ~x[6];
			partial_clause[3][33] 	= partial_clause_prev[3][33] & ~x[5] & ~x[6];
			partial_clause[3][34] 	= partial_clause_prev[3][34] & ~x[2] & ~x[3] & ~x[6];
			partial_clause[3][35] 	= partial_clause_prev[3][35] & ~x[3] & ~x[4] & ~x[5];
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & ~x[5];
			partial_clause[3][38] 	= partial_clause_prev[3][38] & ~x[4] & ~x[6];
			partial_clause[3][39] 	= partial_clause_prev[3][39] & ~x[2] & ~x[4] & ~x[6];
			partial_clause[3][40] 	= partial_clause_prev[3][40] & ~x[6];
			partial_clause[3][41] 	= partial_clause_prev[3][41] & ~x[4] & ~x[6];
			partial_clause[3][42] 	= partial_clause_prev[3][42] & ~x[2] & ~x[6];
			partial_clause[3][43] 	= partial_clause_prev[3][43] & ~x[5];
			partial_clause[3][44] 	= partial_clause_prev[3][44] & ~x[2] & ~x[5];
			partial_clause[3][45] 	= partial_clause_prev[3][45] & ~x[21];
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & ~x[3] & ~x[5];
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & ~x[24];
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & ~x[52];
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & 1'b1;
			partial_clause[3][56] 	= partial_clause_prev[3][56] & ~x[51];
			partial_clause[3][57] 	= partial_clause_prev[3][57] & ~x[52];
			partial_clause[3][58] 	= partial_clause_prev[3][58] & x[5] & ~x[52];
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & ~x[53];
			partial_clause[3][65] 	= partial_clause_prev[3][65] & 1'b1;
			partial_clause[3][66] 	= partial_clause_prev[3][66] & ~x[52];
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & ~x[48];
			partial_clause[3][69] 	= partial_clause_prev[3][69] & ~x[23];
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & ~x[24];
			partial_clause[3][72] 	= partial_clause_prev[3][72] & ~x[47];
			partial_clause[3][73] 	= partial_clause_prev[3][73] & ~x[50] & ~x[52];
			partial_clause[3][74] 	= partial_clause_prev[3][74] & x[5];
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & ~x[40];
			partial_clause[3][78] 	= partial_clause_prev[3][78] & ~x[52];
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & ~x[22];
			partial_clause[3][82] 	= partial_clause_prev[3][82] & ~x[23];
			partial_clause[3][83] 	= partial_clause_prev[3][83] & ~x[52];
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & ~x[23];
			partial_clause[3][87] 	= partial_clause_prev[3][87] & ~x[53];
			partial_clause[3][88] 	= partial_clause_prev[3][88] & x[5] & ~x[51];
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & ~x[42] & ~x[53];
			partial_clause[3][93] 	= partial_clause_prev[3][93] & ~x[25];
			partial_clause[3][94] 	= partial_clause_prev[3][94] & ~x[24] & x[33];
			partial_clause[3][95] 	= partial_clause_prev[3][95] & ~x[50];
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & x[5];
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & ~x[52];
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & ~x[54] & ~x[57];
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & ~x[56];
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & ~x[54];
			partial_clause[4][5] 	= partial_clause_prev[4][5] & ~x[57];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & ~x[56];
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & ~x[14];
			partial_clause[4][14] 	= partial_clause_prev[4][14] & ~x[56];
			partial_clause[4][15] 	= partial_clause_prev[4][15] & ~x[50] & ~x[58];
			partial_clause[4][16] 	= partial_clause_prev[4][16] & ~x[58];
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & ~x[43] & ~x[58];
			partial_clause[4][19] 	= partial_clause_prev[4][19] & ~x[24] & ~x[57];
			partial_clause[4][20] 	= partial_clause_prev[4][20] & ~x[53];
			partial_clause[4][21] 	= partial_clause_prev[4][21] & ~x[58];
			partial_clause[4][22] 	= partial_clause_prev[4][22] & ~x[55];
			partial_clause[4][23] 	= partial_clause_prev[4][23] & ~x[16];
			partial_clause[4][24] 	= partial_clause_prev[4][24] & ~x[15] & ~x[57];
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & ~x[58];
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & ~x[56];
			partial_clause[4][29] 	= partial_clause_prev[4][29] & ~x[25] & ~x[58];
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[57];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & ~x[29] & ~x[51];
			partial_clause[4][35] 	= partial_clause_prev[4][35] & ~x[56];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & ~x[55];
			partial_clause[4][37] 	= partial_clause_prev[4][37] & ~x[56];
			partial_clause[4][38] 	= partial_clause_prev[4][38] & ~x[56];
			partial_clause[4][39] 	= partial_clause_prev[4][39] & ~x[56];
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & ~x[57];
			partial_clause[4][43] 	= partial_clause_prev[4][43] & ~x[30] & ~x[55];
			partial_clause[4][44] 	= partial_clause_prev[4][44] & ~x[31] & ~x[53];
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & ~x[16] & ~x[57];
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & ~x[55] & ~x[58];
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[52] & ~x[57];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & ~x[49];
			partial_clause[4][51] 	= partial_clause_prev[4][51] & ~x[45] & ~x[46];
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & ~x[17];
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & ~x[44];
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & x[57];
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & ~x[50];
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & ~x[47];
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & ~x[22] & ~x[47] & ~x[50];
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & ~x[4];
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & ~x[3] & ~x[4] & ~x[45];
			partial_clause[5][4] 	= partial_clause_prev[5][4] & ~x[15];
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & ~x[2] & ~x[5];
			partial_clause[5][7] 	= partial_clause_prev[5][7] & ~x[3];
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & ~x[3] & ~x[4] & ~x[6];
			partial_clause[5][11] 	= partial_clause_prev[5][11] & ~x[3];
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & ~x[2] & ~x[3];
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & ~x[6];
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & ~x[2] & ~x[3];
			partial_clause[5][19] 	= partial_clause_prev[5][19] & ~x[4];
			partial_clause[5][20] 	= partial_clause_prev[5][20] & ~x[3];
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & ~x[3];
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & ~x[49];
			partial_clause[5][28] 	= partial_clause_prev[5][28] & ~x[33] & ~x[50];
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & ~x[3] & ~x[5];
			partial_clause[5][31] 	= partial_clause_prev[5][31] & ~x[3] & ~x[5];
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & ~x[3];
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & ~x[3];
			partial_clause[5][37] 	= partial_clause_prev[5][37] & ~x[20];
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & ~x[4] & ~x[5];
			partial_clause[5][40] 	= partial_clause_prev[5][40] & ~x[3] & ~x[6];
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & ~x[13];
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & ~x[4] & ~x[6];
			partial_clause[5][49] 	= partial_clause_prev[5][49] & ~x[3];
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & x[34];
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & ~x[44];
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & ~x[54];
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & x[2];
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & x[5];
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & ~x[49];
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & ~x[21];
			partial_clause[5][93] 	= partial_clause_prev[5][93] & ~x[18];
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & x[6];
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & x[31] & x[61] & x[63];
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & x[63];
			partial_clause[6][6] 	= partial_clause_prev[6][6] & x[31];
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & x[60];
			partial_clause[6][9] 	= partial_clause_prev[6][9] & x[60];
			partial_clause[6][10] 	= partial_clause_prev[6][10] & x[60];
			partial_clause[6][11] 	= partial_clause_prev[6][11] & x[31] & ~x[46] & x[61];
			partial_clause[6][12] 	= partial_clause_prev[6][12] & x[2];
			partial_clause[6][13] 	= partial_clause_prev[6][13] & x[60];
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & x[61];
			partial_clause[6][19] 	= partial_clause_prev[6][19] & x[60];
			partial_clause[6][20] 	= partial_clause_prev[6][20] & x[30];
			partial_clause[6][21] 	= partial_clause_prev[6][21] & x[30];
			partial_clause[6][22] 	= partial_clause_prev[6][22] & x[31];
			partial_clause[6][23] 	= partial_clause_prev[6][23] & ~x[17] & x[60];
			partial_clause[6][24] 	= partial_clause_prev[6][24] & x[60];
			partial_clause[6][25] 	= partial_clause_prev[6][25] & ~x[24];
			partial_clause[6][26] 	= partial_clause_prev[6][26] & x[60];
			partial_clause[6][27] 	= partial_clause_prev[6][27] & x[31];
			partial_clause[6][28] 	= partial_clause_prev[6][28] & x[63];
			partial_clause[6][29] 	= partial_clause_prev[6][29] & x[2];
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & x[59];
			partial_clause[6][35] 	= partial_clause_prev[6][35] & x[37];
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & x[31];
			partial_clause[6][39] 	= partial_clause_prev[6][39] & x[63];
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & x[31];
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & x[60];
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & ~x[2];
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & ~x[31];
			partial_clause[6][56] 	= partial_clause_prev[6][56] & ~x[2];
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & ~x[2];
			partial_clause[6][63] 	= partial_clause_prev[6][63] & ~x[1];
			partial_clause[6][64] 	= partial_clause_prev[6][64] & ~x[2];
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & ~x[2];
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & ~x[12];
			partial_clause[6][73] 	= partial_clause_prev[6][73] & ~x[2];
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & ~x[3] & ~x[30];
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & ~x[31];
			partial_clause[6][92] 	= partial_clause_prev[6][92] & ~x[19];
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & ~x[3];
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & ~x[2];
			partial_clause[6][97] 	= partial_clause_prev[6][97] & ~x[31];
			partial_clause[6][98] 	= partial_clause_prev[6][98] & ~x[31];
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & ~x[13] & ~x[57];
			partial_clause[7][1] 	= partial_clause_prev[7][1] & ~x[26];
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & ~x[56];
			partial_clause[7][4] 	= partial_clause_prev[7][4] & ~x[27];
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & ~x[1] & ~x[15] & ~x[27] & ~x[42] & ~x[54];
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & ~x[57];
			partial_clause[7][9] 	= partial_clause_prev[7][9] & ~x[2];
			partial_clause[7][10] 	= partial_clause_prev[7][10] & ~x[28];
			partial_clause[7][11] 	= partial_clause_prev[7][11] & ~x[0] & ~x[26] & ~x[29];
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & ~x[56];
			partial_clause[7][15] 	= partial_clause_prev[7][15] & ~x[54] & ~x[57];
			partial_clause[7][16] 	= partial_clause_prev[7][16] & ~x[2];
			partial_clause[7][17] 	= partial_clause_prev[7][17] & ~x[26];
			partial_clause[7][18] 	= partial_clause_prev[7][18] & ~x[26] & ~x[29];
			partial_clause[7][19] 	= partial_clause_prev[7][19] & ~x[13] & ~x[27];
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & ~x[43] & ~x[55];
			partial_clause[7][22] 	= partial_clause_prev[7][22] & ~x[28];
			partial_clause[7][23] 	= partial_clause_prev[7][23] & ~x[15] & ~x[41];
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & ~x[28];
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & ~x[1] & ~x[2] & ~x[54];
			partial_clause[7][29] 	= partial_clause_prev[7][29] & ~x[56];
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & ~x[27];
			partial_clause[7][32] 	= partial_clause_prev[7][32] & ~x[0] & ~x[56];
			partial_clause[7][33] 	= partial_clause_prev[7][33] & ~x[14];
			partial_clause[7][34] 	= partial_clause_prev[7][34] & ~x[0];
			partial_clause[7][35] 	= partial_clause_prev[7][35] & ~x[29];
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & ~x[19] & ~x[27];
			partial_clause[7][38] 	= partial_clause_prev[7][38] & ~x[26];
			partial_clause[7][39] 	= partial_clause_prev[7][39] & ~x[13];
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & ~x[1];
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & ~x[54];
			partial_clause[7][44] 	= partial_clause_prev[7][44] & ~x[46];
			partial_clause[7][45] 	= partial_clause_prev[7][45] & ~x[1] & ~x[54];
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & ~x[28];
			partial_clause[7][48] 	= partial_clause_prev[7][48] & ~x[26];
			partial_clause[7][49] 	= partial_clause_prev[7][49] & ~x[50];
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & x[38];
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & ~x[46];
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & ~x[49];
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & x[38];
			partial_clause[7][90] 	= partial_clause_prev[7][90] & ~x[19] & x[57];
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & x[3];
			partial_clause[8][1] 	= partial_clause_prev[8][1] & x[3];
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & ~x[47];
			partial_clause[8][5] 	= partial_clause_prev[8][5] & ~x[25];
			partial_clause[8][6] 	= partial_clause_prev[8][6] & x[3] & ~x[23] & ~x[45];
			partial_clause[8][7] 	= partial_clause_prev[8][7] & x[2];
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & x[2];
			partial_clause[8][10] 	= partial_clause_prev[8][10] & x[2];
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & ~x[52];
			partial_clause[8][13] 	= partial_clause_prev[8][13] & x[3] & ~x[24];
			partial_clause[8][14] 	= partial_clause_prev[8][14] & ~x[22];
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & x[3];
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & ~x[16];
			partial_clause[8][19] 	= partial_clause_prev[8][19] & x[2];
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & x[2];
			partial_clause[8][22] 	= partial_clause_prev[8][22] & ~x[25] & x[30];
			partial_clause[8][23] 	= partial_clause_prev[8][23] & ~x[24];
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & ~x[51];
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & x[3] & ~x[52];
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & x[3] & ~x[41];
			partial_clause[8][31] 	= partial_clause_prev[8][31] & x[2];
			partial_clause[8][32] 	= partial_clause_prev[8][32] & x[2];
			partial_clause[8][33] 	= partial_clause_prev[8][33] & x[2] & ~x[43];
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & x[3];
			partial_clause[8][36] 	= partial_clause_prev[8][36] & x[30];
			partial_clause[8][37] 	= partial_clause_prev[8][37] & x[3];
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & ~x[49];
			partial_clause[8][40] 	= partial_clause_prev[8][40] & x[30];
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & x[2] & ~x[20];
			partial_clause[8][43] 	= partial_clause_prev[8][43] & x[2] & ~x[46];
			partial_clause[8][44] 	= partial_clause_prev[8][44] & ~x[16];
			partial_clause[8][45] 	= partial_clause_prev[8][45] & ~x[15];
			partial_clause[8][46] 	= partial_clause_prev[8][46] & x[3];
			partial_clause[8][47] 	= partial_clause_prev[8][47] & x[3];
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & ~x[23];
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & ~x[4] & ~x[20];
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & ~x[1] & ~x[4] & ~x[30];
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & ~x[50];
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & ~x[1] & ~x[2] & ~x[3] & ~x[4];
			partial_clause[8][77] 	= partial_clause_prev[8][77] & ~x[27] & ~x[31] & ~x[57];
			partial_clause[8][78] 	= partial_clause_prev[8][78] & ~x[0] & ~x[2] & ~x[4];
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & ~x[47];
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & 1'b1;
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & ~x[43];
			partial_clause[8][97] 	= partial_clause_prev[8][97] & ~x[51];
			partial_clause[8][98] 	= partial_clause_prev[8][98] & ~x[0] & ~x[28] & ~x[29] & ~x[32];
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & ~x[27] & ~x[58];
			partial_clause[9][1] 	= partial_clause_prev[9][1] & ~x[54] & ~x[57];
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & ~x[42];
			partial_clause[9][4] 	= partial_clause_prev[9][4] & ~x[58];
			partial_clause[9][5] 	= partial_clause_prev[9][5] & ~x[26] & ~x[29];
			partial_clause[9][6] 	= partial_clause_prev[9][6] & ~x[55] & ~x[56] & ~x[58];
			partial_clause[9][7] 	= partial_clause_prev[9][7] & ~x[28] & ~x[31];
			partial_clause[9][8] 	= partial_clause_prev[9][8] & ~x[57];
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & ~x[57] & ~x[58] & ~x[59];
			partial_clause[9][11] 	= partial_clause_prev[9][11] & ~x[55];
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & ~x[30];
			partial_clause[9][14] 	= partial_clause_prev[9][14] & ~x[14] & ~x[49] & ~x[57];
			partial_clause[9][15] 	= partial_clause_prev[9][15] & ~x[56];
			partial_clause[9][16] 	= partial_clause_prev[9][16] & ~x[60];
			partial_clause[9][17] 	= partial_clause_prev[9][17] & ~x[58];
			partial_clause[9][18] 	= partial_clause_prev[9][18] & ~x[12] & ~x[42] & ~x[56];
			partial_clause[9][19] 	= partial_clause_prev[9][19] & ~x[59];
			partial_clause[9][20] 	= partial_clause_prev[9][20] & ~x[56];
			partial_clause[9][21] 	= partial_clause_prev[9][21] & ~x[42] & ~x[57];
			partial_clause[9][22] 	= partial_clause_prev[9][22] & ~x[54];
			partial_clause[9][23] 	= partial_clause_prev[9][23] & ~x[57];
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & ~x[57];
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & ~x[59];
			partial_clause[9][28] 	= partial_clause_prev[9][28] & ~x[56];
			partial_clause[9][29] 	= partial_clause_prev[9][29] & ~x[57];
			partial_clause[9][30] 	= partial_clause_prev[9][30] & ~x[27];
			partial_clause[9][31] 	= partial_clause_prev[9][31] & ~x[41] & ~x[56];
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & ~x[56] & ~x[57];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & ~x[29];
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & ~x[56];
			partial_clause[9][39] 	= partial_clause_prev[9][39] & ~x[28] & ~x[57];
			partial_clause[9][40] 	= partial_clause_prev[9][40] & ~x[57];
			partial_clause[9][41] 	= partial_clause_prev[9][41] & ~x[56];
			partial_clause[9][42] 	= partial_clause_prev[9][42] & ~x[27] & ~x[56];
			partial_clause[9][43] 	= partial_clause_prev[9][43] & ~x[29];
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & ~x[57];
			partial_clause[9][46] 	= partial_clause_prev[9][46] & ~x[55];
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & ~x[56];
			partial_clause[9][49] 	= partial_clause_prev[9][49] & ~x[53];
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & ~x[20];
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & x[57];
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & ~x[49];
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & 1'b1;
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & ~x[46];
			partial_clause[9][75] 	= partial_clause_prev[9][75] & 1'b1;
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & x[56];
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
		end
	end
endmodule


module HCB_9 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & x[22];
			partial_clause[0][1] 	= partial_clause_prev[0][1] & x[21];
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & x[52];
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & ~x[61];
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & 1'b1;
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & x[22];
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & ~x[14];
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & ~x[15];
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & ~x[35];
			partial_clause[0][50] 	= partial_clause_prev[0][50] & ~x[36];
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & ~x[14];
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & ~x[45];
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & ~x[38];
			partial_clause[0][63] 	= partial_clause_prev[0][63] & ~x[13];
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & ~x[11];
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & ~x[41];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & ~x[40];
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & ~x[14];
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & ~x[41];
			partial_clause[0][88] 	= partial_clause_prev[0][88] & 1'b1;
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & 1'b1;
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & ~x[12];
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & 1'b1;
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & ~x[41];
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & ~x[2] & ~x[60];
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & ~x[2];
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & ~x[32];
			partial_clause[1][8] 	= partial_clause_prev[1][8] & ~x[61];
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & ~x[30];
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & ~x[2];
			partial_clause[1][20] 	= partial_clause_prev[1][20] & ~x[46];
			partial_clause[1][21] 	= partial_clause_prev[1][21] & ~x[4];
			partial_clause[1][22] 	= partial_clause_prev[1][22] & ~x[33];
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & ~x[2];
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & ~x[3];
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & ~x[4] & ~x[16];
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & ~x[3];
			partial_clause[1][31] 	= partial_clause_prev[1][31] & ~x[2];
			partial_clause[1][32] 	= partial_clause_prev[1][32] & ~x[30];
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & ~x[3];
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & ~x[2];
			partial_clause[1][41] 	= partial_clause_prev[1][41] & ~x[33];
			partial_clause[1][42] 	= partial_clause_prev[1][42] & ~x[31];
			partial_clause[1][43] 	= partial_clause_prev[1][43] & ~x[2] & ~x[59];
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & ~x[2];
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & ~x[42];
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & ~x[39];
			partial_clause[1][54] 	= partial_clause_prev[1][54] & ~x[13] & ~x[43];
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & ~x[42];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & 1'b1;
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & ~x[38];
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & ~x[36] & ~x[41];
			partial_clause[1][70] 	= partial_clause_prev[1][70] & ~x[38];
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & ~x[37];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & ~x[41];
			partial_clause[1][76] 	= partial_clause_prev[1][76] & ~x[42];
			partial_clause[1][77] 	= partial_clause_prev[1][77] & ~x[9];
			partial_clause[1][78] 	= partial_clause_prev[1][78] & ~x[13];
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & 1'b1;
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & ~x[10];
			partial_clause[1][90] 	= partial_clause_prev[1][90] & ~x[41];
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & ~x[15];
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & ~x[37];
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & 1'b1;
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & ~x[39];
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & ~x[40];
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & 1'b1;
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & ~x[5] & ~x[33] & ~x[37];
			partial_clause[2][51] 	= partial_clause_prev[2][51] & ~x[5] & ~x[31] & ~x[61];
			partial_clause[2][52] 	= partial_clause_prev[2][52] & ~x[7] & ~x[20] & ~x[60];
			partial_clause[2][53] 	= partial_clause_prev[2][53] & ~x[5] & ~x[7];
			partial_clause[2][54] 	= partial_clause_prev[2][54] & ~x[4] & ~x[61];
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & ~x[6];
			partial_clause[2][57] 	= partial_clause_prev[2][57] & ~x[14] & ~x[33];
			partial_clause[2][58] 	= partial_clause_prev[2][58] & ~x[5];
			partial_clause[2][59] 	= partial_clause_prev[2][59] & ~x[5] & ~x[8] & ~x[60];
			partial_clause[2][60] 	= partial_clause_prev[2][60] & ~x[5] & ~x[19] & ~x[60];
			partial_clause[2][61] 	= partial_clause_prev[2][61] & ~x[7] & ~x[31] & ~x[35] & ~x[44];
			partial_clause[2][62] 	= partial_clause_prev[2][62] & ~x[35] & ~x[60];
			partial_clause[2][63] 	= partial_clause_prev[2][63] & ~x[33] & ~x[62] & ~x[63];
			partial_clause[2][64] 	= partial_clause_prev[2][64] & ~x[6];
			partial_clause[2][65] 	= partial_clause_prev[2][65] & ~x[5] & ~x[35];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & ~x[32] & ~x[61];
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & ~x[7];
			partial_clause[2][70] 	= partial_clause_prev[2][70] & ~x[5] & ~x[6] & ~x[60];
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & ~x[6] & ~x[34];
			partial_clause[2][73] 	= partial_clause_prev[2][73] & ~x[4];
			partial_clause[2][74] 	= partial_clause_prev[2][74] & ~x[34] & ~x[63];
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & ~x[7] & ~x[62] & ~x[63];
			partial_clause[2][77] 	= partial_clause_prev[2][77] & ~x[7];
			partial_clause[2][78] 	= partial_clause_prev[2][78] & ~x[60];
			partial_clause[2][79] 	= partial_clause_prev[2][79] & ~x[6] & ~x[7];
			partial_clause[2][80] 	= partial_clause_prev[2][80] & ~x[33];
			partial_clause[2][81] 	= partial_clause_prev[2][81] & ~x[32];
			partial_clause[2][82] 	= partial_clause_prev[2][82] & ~x[4] & ~x[59];
			partial_clause[2][83] 	= partial_clause_prev[2][83] & ~x[4] & ~x[59];
			partial_clause[2][84] 	= partial_clause_prev[2][84] & ~x[32] & ~x[33] & ~x[59];
			partial_clause[2][85] 	= partial_clause_prev[2][85] & ~x[6] & ~x[34];
			partial_clause[2][86] 	= partial_clause_prev[2][86] & ~x[6];
			partial_clause[2][87] 	= partial_clause_prev[2][87] & ~x[44];
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & ~x[39];
			partial_clause[2][90] 	= partial_clause_prev[2][90] & ~x[62];
			partial_clause[2][91] 	= partial_clause_prev[2][91] & ~x[35];
			partial_clause[2][92] 	= partial_clause_prev[2][92] & ~x[35];
			partial_clause[2][93] 	= partial_clause_prev[2][93] & ~x[7];
			partial_clause[2][94] 	= partial_clause_prev[2][94] & ~x[7] & ~x[33];
			partial_clause[2][95] 	= partial_clause_prev[2][95] & ~x[5];
			partial_clause[2][96] 	= partial_clause_prev[2][96] & ~x[35];
			partial_clause[2][97] 	= partial_clause_prev[2][97] & ~x[8] & ~x[17] & ~x[35];
			partial_clause[2][98] 	= partial_clause_prev[2][98] & ~x[7];
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & ~x[12];
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & ~x[35];
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & ~x[13];
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & ~x[7] & ~x[41];
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & ~x[11];
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & ~x[63];
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & ~x[40];
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & ~x[45];
			partial_clause[3][52] 	= partial_clause_prev[3][52] & ~x[43] & ~x[46];
			partial_clause[3][53] 	= partial_clause_prev[3][53] & ~x[43];
			partial_clause[3][54] 	= partial_clause_prev[3][54] & ~x[16] & ~x[46];
			partial_clause[3][55] 	= partial_clause_prev[3][55] & ~x[41];
			partial_clause[3][56] 	= partial_clause_prev[3][56] & ~x[44];
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & ~x[48] & ~x[49] & ~x[58];
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & ~x[16];
			partial_clause[3][64] 	= partial_clause_prev[3][64] & ~x[18];
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[16];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & ~x[42];
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & ~x[59];
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & ~x[9] & ~x[13] & ~x[47];
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & ~x[45];
			partial_clause[3][76] 	= partial_clause_prev[3][76] & ~x[17];
			partial_clause[3][77] 	= partial_clause_prev[3][77] & ~x[38];
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & ~x[16];
			partial_clause[3][80] 	= partial_clause_prev[3][80] & ~x[44];
			partial_clause[3][81] 	= partial_clause_prev[3][81] & ~x[42];
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & ~x[16] & ~x[17] & ~x[45];
			partial_clause[3][84] 	= partial_clause_prev[3][84] & ~x[17] & ~x[47];
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & ~x[41];
			partial_clause[3][87] 	= partial_clause_prev[3][87] & ~x[8];
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & ~x[19];
			partial_clause[3][90] 	= partial_clause_prev[3][90] & ~x[14] & ~x[42];
			partial_clause[3][91] 	= partial_clause_prev[3][91] & ~x[17] & ~x[46];
			partial_clause[3][92] 	= partial_clause_prev[3][92] & ~x[16];
			partial_clause[3][93] 	= partial_clause_prev[3][93] & ~x[48];
			partial_clause[3][94] 	= partial_clause_prev[3][94] & ~x[16];
			partial_clause[3][95] 	= partial_clause_prev[3][95] & ~x[15];
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & ~x[17] & ~x[45];
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & ~x[46];
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & ~x[20];
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & ~x[48];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & ~x[17];
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & ~x[19];
			partial_clause[4][11] 	= partial_clause_prev[4][11] & ~x[20];
			partial_clause[4][12] 	= partial_clause_prev[4][12] & ~x[48];
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & ~x[16];
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & ~x[21];
			partial_clause[4][17] 	= partial_clause_prev[4][17] & ~x[40];
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & ~x[19];
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & ~x[20];
			partial_clause[4][24] 	= partial_clause_prev[4][24] & ~x[49];
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & ~x[49];
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & ~x[48];
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & 1'b1;
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & ~x[47];
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & ~x[20];
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & ~x[19] & ~x[40];
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & ~x[11] & ~x[19] & ~x[21];
			partial_clause[4][45] 	= partial_clause_prev[4][45] & ~x[19];
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & ~x[19];
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & 1'b1;
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & x[52];
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & 1'b1;
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & x[51] & x[54];
			partial_clause[4][69] 	= partial_clause_prev[4][69] & x[23];
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & ~x[14] & ~x[42];
			partial_clause[4][73] 	= partial_clause_prev[4][73] & ~x[13] & x[52];
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & ~x[13];
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & ~x[42];
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & ~x[10];
			partial_clause[4][80] 	= partial_clause_prev[4][80] & x[21];
			partial_clause[4][81] 	= partial_clause_prev[4][81] & ~x[14];
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & x[19];
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & x[21];
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & x[23] & ~x[42];
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & ~x[13];
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & x[21] & ~x[41];
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & ~x[11];
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & ~x[9];
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & ~x[40];
			partial_clause[5][52] 	= partial_clause_prev[5][52] & ~x[11] & ~x[59];
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & ~x[63];
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & ~x[57];
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & ~x[44];
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & ~x[37];
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & ~x[15];
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & ~x[37];
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & ~x[38];
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & ~x[59];
			partial_clause[6][1] 	= partial_clause_prev[6][1] & ~x[12];
			partial_clause[6][2] 	= partial_clause_prev[6][2] & ~x[35];
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & ~x[48];
			partial_clause[6][5] 	= partial_clause_prev[6][5] & ~x[18] & ~x[48];
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & ~x[47] & ~x[48] & ~x[49];
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & ~x[48];
			partial_clause[6][11] 	= partial_clause_prev[6][11] & ~x[18];
			partial_clause[6][12] 	= partial_clause_prev[6][12] & ~x[46];
			partial_clause[6][13] 	= partial_clause_prev[6][13] & ~x[49] & ~x[62];
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & ~x[9];
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & ~x[18] & ~x[40];
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & ~x[47];
			partial_clause[6][21] 	= partial_clause_prev[6][21] & ~x[46];
			partial_clause[6][22] 	= partial_clause_prev[6][22] & ~x[45] & ~x[49];
			partial_clause[6][23] 	= partial_clause_prev[6][23] & ~x[19];
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & ~x[8] & ~x[49];
			partial_clause[6][27] 	= partial_clause_prev[6][27] & ~x[9];
			partial_clause[6][28] 	= partial_clause_prev[6][28] & ~x[33];
			partial_clause[6][29] 	= partial_clause_prev[6][29] & ~x[34];
			partial_clause[6][30] 	= partial_clause_prev[6][30] & ~x[7] & ~x[60];
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & ~x[8];
			partial_clause[6][34] 	= partial_clause_prev[6][34] & ~x[48];
			partial_clause[6][35] 	= partial_clause_prev[6][35] & ~x[35];
			partial_clause[6][36] 	= partial_clause_prev[6][36] & ~x[46];
			partial_clause[6][37] 	= partial_clause_prev[6][37] & ~x[36] & ~x[49];
			partial_clause[6][38] 	= partial_clause_prev[6][38] & ~x[19];
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & ~x[47];
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & ~x[7] & ~x[59];
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & ~x[15] & ~x[61];
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & ~x[42];
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & ~x[14];
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & ~x[12];
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & ~x[12];
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & ~x[18];
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & ~x[34];
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & ~x[19];
			partial_clause[7][10] 	= partial_clause_prev[7][10] & ~x[4] & ~x[5];
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & ~x[20];
			partial_clause[7][13] 	= partial_clause_prev[7][13] & ~x[5];
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & ~x[19];
			partial_clause[7][16] 	= partial_clause_prev[7][16] & ~x[5] & ~x[19] & ~x[45];
			partial_clause[7][17] 	= partial_clause_prev[7][17] & ~x[33];
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & ~x[32];
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & ~x[18];
			partial_clause[7][22] 	= partial_clause_prev[7][22] & ~x[18];
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & ~x[36];
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & ~x[5] & ~x[20];
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & ~x[19];
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & ~x[19];
			partial_clause[7][37] 	= partial_clause_prev[7][37] & ~x[19];
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & ~x[44];
			partial_clause[7][41] 	= partial_clause_prev[7][41] & ~x[19] & ~x[33];
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & ~x[15];
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & 1'b1;
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & ~x[12];
			partial_clause[7][57] 	= partial_clause_prev[7][57] & ~x[12];
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & 1'b1;
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & x[20];
			partial_clause[7][78] 	= partial_clause_prev[7][78] & 1'b1;
			partial_clause[7][79] 	= partial_clause_prev[7][79] & ~x[42];
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & 1'b1;
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & 1'b1;
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & ~x[14];
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & ~x[40];
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & 1'b1;
			partial_clause[8][25] 	= partial_clause_prev[8][25] & ~x[63];
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & ~x[38];
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & ~x[13];
			partial_clause[8][48] 	= partial_clause_prev[8][48] & ~x[34] & ~x[44];
			partial_clause[8][49] 	= partial_clause_prev[8][49] & x[53];
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & ~x[41] & ~x[42];
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & ~x[12];
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & ~x[51] & ~x[58];
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & ~x[62];
			partial_clause[8][58] 	= partial_clause_prev[8][58] & ~x[7];
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & ~x[35] & ~x[47];
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & ~x[22] & ~x[47] & ~x[49];
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & ~x[37];
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & ~x[9];
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & ~x[40];
			partial_clause[8][85] 	= partial_clause_prev[8][85] & ~x[50];
			partial_clause[8][86] 	= partial_clause_prev[8][86] & 1'b1;
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & 1'b1;
			partial_clause[8][90] 	= partial_clause_prev[8][90] & ~x[39];
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & ~x[51] & ~x[58];
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & ~x[46] & ~x[47] & ~x[48];
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & ~x[20] & ~x[38] & ~x[48];
			partial_clause[9][2] 	= partial_clause_prev[9][2] & ~x[20];
			partial_clause[9][3] 	= partial_clause_prev[9][3] & ~x[22];
			partial_clause[9][4] 	= partial_clause_prev[9][4] & ~x[47];
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & ~x[48];
			partial_clause[9][7] 	= partial_clause_prev[9][7] & ~x[19] & ~x[21];
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & ~x[50];
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & ~x[19];
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & ~x[21];
			partial_clause[9][16] 	= partial_clause_prev[9][16] & ~x[22];
			partial_clause[9][17] 	= partial_clause_prev[9][17] & ~x[47];
			partial_clause[9][18] 	= partial_clause_prev[9][18] & ~x[44];
			partial_clause[9][19] 	= partial_clause_prev[9][19] & ~x[20] & ~x[23];
			partial_clause[9][20] 	= partial_clause_prev[9][20] & ~x[18];
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & ~x[22] & ~x[47] & ~x[62];
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & ~x[48];
			partial_clause[9][25] 	= partial_clause_prev[9][25] & ~x[20];
			partial_clause[9][26] 	= partial_clause_prev[9][26] & ~x[17];
			partial_clause[9][27] 	= partial_clause_prev[9][27] & ~x[48] & ~x[50];
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & ~x[47];
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & ~x[20];
			partial_clause[9][33] 	= partial_clause_prev[9][33] & ~x[22] & ~x[49];
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & ~x[20];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & ~x[50];
			partial_clause[9][39] 	= partial_clause_prev[9][39] & ~x[47];
			partial_clause[9][40] 	= partial_clause_prev[9][40] & ~x[18];
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & ~x[19];
			partial_clause[9][44] 	= partial_clause_prev[9][44] & ~x[19];
			partial_clause[9][45] 	= partial_clause_prev[9][45] & ~x[20];
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & ~x[47];
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & ~x[12];
			partial_clause[9][52] 	= partial_clause_prev[9][52] & ~x[12];
			partial_clause[9][53] 	= partial_clause_prev[9][53] & x[50];
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & ~x[11] & x[22] & ~x[39];
			partial_clause[9][56] 	= partial_clause_prev[9][56] & 1'b1;
			partial_clause[9][57] 	= partial_clause_prev[9][57] & x[22];
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & x[23];
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & ~x[63];
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & x[22];
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & x[51];
			partial_clause[9][73] 	= partial_clause_prev[9][73] & x[21];
			partial_clause[9][74] 	= partial_clause_prev[9][74] & x[21];
			partial_clause[9][75] 	= partial_clause_prev[9][75] & x[23];
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & x[26];
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & x[24];
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & x[49];
			partial_clause[9][92] 	= partial_clause_prev[9][92] & ~x[11];
			partial_clause[9][93] 	= partial_clause_prev[9][93] & x[20];
			partial_clause[9][94] 	= partial_clause_prev[9][94] & ~x[37];
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
		end
	end
endmodule


module HCB_10 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & ~x[35];
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & ~x[3];
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & ~x[36];
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & ~x[37];
			partial_clause[0][14] 	= partial_clause_prev[0][14] & ~x[3];
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & ~x[50];
			partial_clause[0][22] 	= partial_clause_prev[0][22] & ~x[8] & ~x[35];
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & ~x[26] & ~x[35];
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & ~x[32];
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & 1'b1;
			partial_clause[0][30] 	= partial_clause_prev[0][30] & x[16];
			partial_clause[0][31] 	= partial_clause_prev[0][31] & ~x[25];
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & ~x[5];
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & ~x[30];
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & 1'b1;
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & ~x[60];
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & ~x[53];
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & ~x[7];
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & 1'b1;
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & ~x[3] & ~x[60];
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & ~x[62];
			partial_clause[0][65] 	= partial_clause_prev[0][65] & ~x[27];
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & ~x[61];
			partial_clause[0][69] 	= partial_clause_prev[0][69] & ~x[34];
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & 1'b1;
			partial_clause[0][73] 	= partial_clause_prev[0][73] & ~x[31];
			partial_clause[0][74] 	= partial_clause_prev[0][74] & ~x[0];
			partial_clause[0][75] 	= partial_clause_prev[0][75] & ~x[60];
			partial_clause[0][76] 	= partial_clause_prev[0][76] & ~x[36];
			partial_clause[0][77] 	= partial_clause_prev[0][77] & ~x[53];
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & ~x[35];
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & ~x[8];
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & ~x[5] & ~x[28];
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & 1'b1;
			partial_clause[0][91] 	= partial_clause_prev[0][91] & ~x[4] & ~x[5];
			partial_clause[0][92] 	= partial_clause_prev[0][92] & ~x[61];
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & ~x[33];
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & ~x[33];
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & ~x[61];
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & ~x[26];
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & ~x[22];
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & ~x[54];
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & ~x[59];
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & ~x[0] & ~x[30] & ~x[31];
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & ~x[3] & ~x[5];
			partial_clause[1][54] 	= partial_clause_prev[1][54] & ~x[36];
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & ~x[63];
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & ~x[8];
			partial_clause[1][59] 	= partial_clause_prev[1][59] & ~x[3] & ~x[37];
			partial_clause[1][60] 	= partial_clause_prev[1][60] & ~x[29];
			partial_clause[1][61] 	= partial_clause_prev[1][61] & 1'b1;
			partial_clause[1][62] 	= partial_clause_prev[1][62] & 1'b1;
			partial_clause[1][63] 	= partial_clause_prev[1][63] & ~x[37];
			partial_clause[1][64] 	= partial_clause_prev[1][64] & ~x[0];
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & ~x[60];
			partial_clause[1][67] 	= partial_clause_prev[1][67] & ~x[6] & ~x[63];
			partial_clause[1][68] 	= partial_clause_prev[1][68] & 1'b1;
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & 1'b1;
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & 1'b1;
			partial_clause[1][74] 	= partial_clause_prev[1][74] & 1'b1;
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & ~x[32];
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & ~x[55];
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & ~x[6] & ~x[32];
			partial_clause[1][88] 	= partial_clause_prev[1][88] & ~x[6];
			partial_clause[1][89] 	= partial_clause_prev[1][89] & ~x[29] & ~x[33];
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & 1'b1;
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & ~x[28];
			partial_clause[1][96] 	= partial_clause_prev[1][96] & ~x[31];
			partial_clause[1][97] 	= partial_clause_prev[1][97] & 1'b1;
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & ~x[56];
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & ~x[16] & ~x[47];
			partial_clause[2][2] 	= partial_clause_prev[2][2] & ~x[47];
			partial_clause[2][3] 	= partial_clause_prev[2][3] & ~x[44];
			partial_clause[2][4] 	= partial_clause_prev[2][4] & ~x[44] & ~x[46];
			partial_clause[2][5] 	= partial_clause_prev[2][5] & ~x[44] & ~x[46];
			partial_clause[2][6] 	= partial_clause_prev[2][6] & ~x[5] & ~x[35] & ~x[44];
			partial_clause[2][7] 	= partial_clause_prev[2][7] & ~x[35] & ~x[44];
			partial_clause[2][8] 	= partial_clause_prev[2][8] & ~x[43];
			partial_clause[2][9] 	= partial_clause_prev[2][9] & ~x[44] & ~x[57];
			partial_clause[2][10] 	= partial_clause_prev[2][10] & ~x[44];
			partial_clause[2][11] 	= partial_clause_prev[2][11] & ~x[41] & ~x[43] & ~x[48];
			partial_clause[2][12] 	= partial_clause_prev[2][12] & ~x[44];
			partial_clause[2][13] 	= partial_clause_prev[2][13] & ~x[43] & ~x[55];
			partial_clause[2][14] 	= partial_clause_prev[2][14] & ~x[38] & ~x[43] & ~x[45];
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & ~x[42];
			partial_clause[2][17] 	= partial_clause_prev[2][17] & ~x[40] & ~x[43] & ~x[46];
			partial_clause[2][18] 	= partial_clause_prev[2][18] & ~x[42];
			partial_clause[2][19] 	= partial_clause_prev[2][19] & ~x[42] & ~x[43] & ~x[46];
			partial_clause[2][20] 	= partial_clause_prev[2][20] & ~x[40] & ~x[41] & ~x[43] & ~x[46];
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & ~x[44];
			partial_clause[2][23] 	= partial_clause_prev[2][23] & ~x[18] & ~x[42] & ~x[48];
			partial_clause[2][24] 	= partial_clause_prev[2][24] & ~x[18];
			partial_clause[2][25] 	= partial_clause_prev[2][25] & ~x[43];
			partial_clause[2][26] 	= partial_clause_prev[2][26] & ~x[44];
			partial_clause[2][27] 	= partial_clause_prev[2][27] & ~x[40] & ~x[41] & ~x[45];
			partial_clause[2][28] 	= partial_clause_prev[2][28] & ~x[41] & ~x[45];
			partial_clause[2][29] 	= partial_clause_prev[2][29] & ~x[44];
			partial_clause[2][30] 	= partial_clause_prev[2][30] & ~x[15] & ~x[44];
			partial_clause[2][31] 	= partial_clause_prev[2][31] & ~x[42] & ~x[43];
			partial_clause[2][32] 	= partial_clause_prev[2][32] & ~x[46];
			partial_clause[2][33] 	= partial_clause_prev[2][33] & ~x[16] & ~x[46];
			partial_clause[2][34] 	= partial_clause_prev[2][34] & ~x[42] & ~x[53];
			partial_clause[2][35] 	= partial_clause_prev[2][35] & ~x[31] & ~x[42];
			partial_clause[2][36] 	= partial_clause_prev[2][36] & ~x[18] & ~x[36] & ~x[44] & ~x[52];
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & ~x[42] & ~x[44] & ~x[47];
			partial_clause[2][39] 	= partial_clause_prev[2][39] & ~x[43];
			partial_clause[2][40] 	= partial_clause_prev[2][40] & ~x[39] & ~x[42];
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & ~x[17] & ~x[48] & ~x[55] & ~x[56];
			partial_clause[2][43] 	= partial_clause_prev[2][43] & ~x[44];
			partial_clause[2][44] 	= partial_clause_prev[2][44] & ~x[41] & ~x[47];
			partial_clause[2][45] 	= partial_clause_prev[2][45] & ~x[18] & ~x[43];
			partial_clause[2][46] 	= partial_clause_prev[2][46] & ~x[42] & ~x[47];
			partial_clause[2][47] 	= partial_clause_prev[2][47] & ~x[18] & ~x[42];
			partial_clause[2][48] 	= partial_clause_prev[2][48] & ~x[18] & ~x[39] & ~x[42] & ~x[43] & ~x[49];
			partial_clause[2][49] 	= partial_clause_prev[2][49] & ~x[40] & ~x[45];
			partial_clause[2][50] 	= partial_clause_prev[2][50] & ~x[25];
			partial_clause[2][51] 	= partial_clause_prev[2][51] & ~x[30];
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & ~x[2] & ~x[58];
			partial_clause[2][59] 	= partial_clause_prev[2][59] & ~x[54];
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & ~x[1];
			partial_clause[2][65] 	= partial_clause_prev[2][65] & ~x[25];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & ~x[34];
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & ~x[25];
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & ~x[3];
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & ~x[2] & ~x[60];
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & ~x[31];
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & ~x[52];
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & ~x[30];
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & 1'b1;
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & ~x[61];
			partial_clause[3][26] 	= partial_clause_prev[3][26] & ~x[5];
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & ~x[33] & ~x[55];
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & ~x[52];
			partial_clause[3][45] 	= partial_clause_prev[3][45] & ~x[4] & ~x[50];
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & ~x[57];
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & ~x[11];
			partial_clause[3][51] 	= partial_clause_prev[3][51] & ~x[39];
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & ~x[7] & ~x[9] & ~x[36];
			partial_clause[3][55] 	= partial_clause_prev[3][55] & ~x[9];
			partial_clause[3][56] 	= partial_clause_prev[3][56] & ~x[8] & ~x[57];
			partial_clause[3][57] 	= partial_clause_prev[3][57] & ~x[32] & ~x[37];
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & ~x[12];
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & ~x[39];
			partial_clause[3][62] 	= partial_clause_prev[3][62] & ~x[32];
			partial_clause[3][63] 	= partial_clause_prev[3][63] & 1'b1;
			partial_clause[3][64] 	= partial_clause_prev[3][64] & ~x[40];
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[10];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & ~x[10];
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & ~x[1];
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & ~x[38] & ~x[62];
			partial_clause[3][71] 	= partial_clause_prev[3][71] & ~x[9];
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & ~x[11];
			partial_clause[3][76] 	= partial_clause_prev[3][76] & ~x[9] & ~x[11];
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & ~x[9];
			partial_clause[3][79] 	= partial_clause_prev[3][79] & ~x[6] & ~x[9] & ~x[39];
			partial_clause[3][80] 	= partial_clause_prev[3][80] & ~x[2] & ~x[11];
			partial_clause[3][81] 	= partial_clause_prev[3][81] & ~x[37] & ~x[63];
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & ~x[30];
			partial_clause[3][84] 	= partial_clause_prev[3][84] & ~x[4] & ~x[37];
			partial_clause[3][85] 	= partial_clause_prev[3][85] & ~x[2] & ~x[6] & ~x[9];
			partial_clause[3][86] 	= partial_clause_prev[3][86] & ~x[11];
			partial_clause[3][87] 	= partial_clause_prev[3][87] & ~x[10];
			partial_clause[3][88] 	= partial_clause_prev[3][88] & ~x[9] & ~x[30] & ~x[37];
			partial_clause[3][89] 	= partial_clause_prev[3][89] & ~x[9] & ~x[11];
			partial_clause[3][90] 	= partial_clause_prev[3][90] & ~x[32];
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & ~x[11];
			partial_clause[3][93] 	= partial_clause_prev[3][93] & ~x[12] & ~x[39];
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & ~x[38];
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & ~x[5];
			partial_clause[4][7] 	= partial_clause_prev[4][7] & 1'b1;
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & ~x[36];
			partial_clause[4][11] 	= partial_clause_prev[4][11] & ~x[0] & ~x[58];
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & ~x[10];
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & ~x[62];
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & 1'b1;
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[0];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & ~x[9];
			partial_clause[4][40] 	= partial_clause_prev[4][40] & ~x[12];
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & ~x[32];
			partial_clause[4][43] 	= partial_clause_prev[4][43] & ~x[3];
			partial_clause[4][44] 	= partial_clause_prev[4][44] & ~x[39];
			partial_clause[4][45] 	= partial_clause_prev[4][45] & ~x[40];
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[31];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & ~x[4];
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & ~x[56];
			partial_clause[4][54] 	= partial_clause_prev[4][54] & ~x[29];
			partial_clause[4][55] 	= partial_clause_prev[4][55] & ~x[56];
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & 1'b1;
			partial_clause[4][59] 	= partial_clause_prev[4][59] & ~x[7];
			partial_clause[4][60] 	= partial_clause_prev[4][60] & ~x[30] & ~x[32] & ~x[61];
			partial_clause[4][61] 	= partial_clause_prev[4][61] & 1'b1;
			partial_clause[4][62] 	= partial_clause_prev[4][62] & ~x[6];
			partial_clause[4][63] 	= partial_clause_prev[4][63] & ~x[29];
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & ~x[22];
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & ~x[52] & ~x[53];
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & ~x[33];
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & ~x[63];
			partial_clause[4][74] 	= partial_clause_prev[4][74] & ~x[3];
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & 1'b1;
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & ~x[25] & ~x[32] & ~x[51];
			partial_clause[4][79] 	= partial_clause_prev[4][79] & ~x[0] & ~x[59];
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & ~x[32] & ~x[56];
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & ~x[63];
			partial_clause[4][85] 	= partial_clause_prev[4][85] & ~x[58];
			partial_clause[4][86] 	= partial_clause_prev[4][86] & ~x[56] & ~x[63];
			partial_clause[4][87] 	= partial_clause_prev[4][87] & ~x[37] & ~x[58];
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & ~x[59];
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & ~x[52] & ~x[57];
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & ~x[62];
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & 1'b1;
			partial_clause[5][9] 	= partial_clause_prev[5][9] & ~x[31];
			partial_clause[5][10] 	= partial_clause_prev[5][10] & ~x[4];
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & ~x[29];
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & ~x[37] & ~x[60];
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & ~x[31];
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & ~x[61];
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & ~x[8];
			partial_clause[5][55] 	= partial_clause_prev[5][55] & ~x[4];
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & ~x[56] & ~x[57];
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & ~x[3];
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & 1'b1;
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & ~x[31];
			partial_clause[5][71] 	= partial_clause_prev[5][71] & ~x[56];
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & 1'b1;
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & ~x[31];
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & ~x[37];
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & ~x[58];
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & ~x[30];
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & ~x[7];
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & ~x[57];
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & ~x[12] & ~x[19];
			partial_clause[6][1] 	= partial_clause_prev[6][1] & ~x[13] & ~x[16] & ~x[20];
			partial_clause[6][2] 	= partial_clause_prev[6][2] & ~x[10] & ~x[14] & ~x[16] & ~x[19] & ~x[49];
			partial_clause[6][3] 	= partial_clause_prev[6][3] & ~x[15] & ~x[19] & ~x[20] & ~x[50];
			partial_clause[6][4] 	= partial_clause_prev[6][4] & ~x[14] & ~x[17] & ~x[18] & ~x[19] & ~x[32];
			partial_clause[6][5] 	= partial_clause_prev[6][5] & ~x[16] & ~x[18] & ~x[20];
			partial_clause[6][6] 	= partial_clause_prev[6][6] & ~x[14] & ~x[21];
			partial_clause[6][7] 	= partial_clause_prev[6][7] & ~x[16] & ~x[19];
			partial_clause[6][8] 	= partial_clause_prev[6][8] & ~x[15] & ~x[47];
			partial_clause[6][9] 	= partial_clause_prev[6][9] & ~x[16] & ~x[18] & ~x[22] & ~x[51];
			partial_clause[6][10] 	= partial_clause_prev[6][10] & ~x[17];
			partial_clause[6][11] 	= partial_clause_prev[6][11] & ~x[16] & ~x[20];
			partial_clause[6][12] 	= partial_clause_prev[6][12] & ~x[13] & ~x[17];
			partial_clause[6][13] 	= partial_clause_prev[6][13] & ~x[16] & ~x[17];
			partial_clause[6][14] 	= partial_clause_prev[6][14] & ~x[18];
			partial_clause[6][15] 	= partial_clause_prev[6][15] & ~x[14] & ~x[19];
			partial_clause[6][16] 	= partial_clause_prev[6][16] & ~x[16] & ~x[17];
			partial_clause[6][17] 	= partial_clause_prev[6][17] & ~x[17] & ~x[19] & ~x[53];
			partial_clause[6][18] 	= partial_clause_prev[6][18] & ~x[45];
			partial_clause[6][19] 	= partial_clause_prev[6][19] & ~x[14] & ~x[17];
			partial_clause[6][20] 	= partial_clause_prev[6][20] & ~x[19] & ~x[25];
			partial_clause[6][21] 	= partial_clause_prev[6][21] & ~x[47];
			partial_clause[6][22] 	= partial_clause_prev[6][22] & ~x[13] & ~x[45];
			partial_clause[6][23] 	= partial_clause_prev[6][23] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[21] & ~x[22];
			partial_clause[6][24] 	= partial_clause_prev[6][24] & ~x[13] & ~x[20] & ~x[43];
			partial_clause[6][25] 	= partial_clause_prev[6][25] & ~x[15];
			partial_clause[6][26] 	= partial_clause_prev[6][26] & ~x[16];
			partial_clause[6][27] 	= partial_clause_prev[6][27] & ~x[13] & ~x[15];
			partial_clause[6][28] 	= partial_clause_prev[6][28] & ~x[13] & ~x[15] & ~x[44] & ~x[45];
			partial_clause[6][29] 	= partial_clause_prev[6][29] & ~x[16] & ~x[20] & ~x[23];
			partial_clause[6][30] 	= partial_clause_prev[6][30] & ~x[14] & ~x[18] & ~x[21];
			partial_clause[6][31] 	= partial_clause_prev[6][31] & ~x[18] & ~x[20] & ~x[45];
			partial_clause[6][32] 	= partial_clause_prev[6][32] & ~x[12] & ~x[18] & ~x[20] & ~x[21] & ~x[43];
			partial_clause[6][33] 	= partial_clause_prev[6][33] & ~x[14] & ~x[16] & ~x[17] & ~x[47];
			partial_clause[6][34] 	= partial_clause_prev[6][34] & ~x[14];
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & ~x[8];
			partial_clause[6][37] 	= partial_clause_prev[6][37] & ~x[16];
			partial_clause[6][38] 	= partial_clause_prev[6][38] & ~x[14] & ~x[17];
			partial_clause[6][39] 	= partial_clause_prev[6][39] & ~x[23];
			partial_clause[6][40] 	= partial_clause_prev[6][40] & ~x[17] & ~x[21] & ~x[38] & ~x[42] & ~x[59];
			partial_clause[6][41] 	= partial_clause_prev[6][41] & ~x[15] & ~x[16] & ~x[18] & ~x[19];
			partial_clause[6][42] 	= partial_clause_prev[6][42] & ~x[25];
			partial_clause[6][43] 	= partial_clause_prev[6][43] & ~x[17] & ~x[18] & ~x[23] & ~x[48];
			partial_clause[6][44] 	= partial_clause_prev[6][44] & ~x[15] & ~x[44];
			partial_clause[6][45] 	= partial_clause_prev[6][45] & ~x[15] & ~x[19];
			partial_clause[6][46] 	= partial_clause_prev[6][46] & ~x[14] & ~x[15] & ~x[19];
			partial_clause[6][47] 	= partial_clause_prev[6][47] & ~x[16] & ~x[19];
			partial_clause[6][48] 	= partial_clause_prev[6][48] & ~x[12] & ~x[18];
			partial_clause[6][49] 	= partial_clause_prev[6][49] & ~x[18] & ~x[19];
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & ~x[30];
			partial_clause[6][53] 	= partial_clause_prev[6][53] & ~x[63];
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & ~x[3];
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & ~x[6];
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & x[17] & ~x[29];
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & ~x[5];
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & ~x[63];
			partial_clause[6][71] 	= partial_clause_prev[6][71] & ~x[0];
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & ~x[32];
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & x[17] & ~x[54];
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & ~x[29];
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & x[15] & ~x[32];
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & 1'b1;
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & ~x[33];
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & x[18];
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & 1'b1;
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & ~x[4];
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & ~x[28];
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & ~x[26];
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & ~x[62];
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & ~x[28];
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & 1'b1;
			partial_clause[7][39] 	= partial_clause_prev[7][39] & ~x[61];
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & ~x[8];
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & ~x[6];
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & ~x[39];
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & 1'b1;
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & ~x[39];
			partial_clause[7][58] 	= partial_clause_prev[7][58] & 1'b1;
			partial_clause[7][59] 	= partial_clause_prev[7][59] & ~x[2] & ~x[39];
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & ~x[38];
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & ~x[37];
			partial_clause[7][65] 	= partial_clause_prev[7][65] & ~x[38];
			partial_clause[7][66] 	= partial_clause_prev[7][66] & 1'b1;
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & ~x[40];
			partial_clause[7][70] 	= partial_clause_prev[7][70] & ~x[38] & ~x[53];
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & ~x[38] & ~x[39] & ~x[41];
			partial_clause[7][73] 	= partial_clause_prev[7][73] & ~x[36] & ~x[37] & ~x[58];
			partial_clause[7][74] 	= partial_clause_prev[7][74] & ~x[2] & ~x[39];
			partial_clause[7][75] 	= partial_clause_prev[7][75] & ~x[55];
			partial_clause[7][76] 	= partial_clause_prev[7][76] & ~x[63];
			partial_clause[7][77] 	= partial_clause_prev[7][77] & ~x[39];
			partial_clause[7][78] 	= partial_clause_prev[7][78] & ~x[39];
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & ~x[38];
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & 1'b1;
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & ~x[37];
			partial_clause[7][88] 	= partial_clause_prev[7][88] & ~x[38] & ~x[40];
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & 1'b1;
			partial_clause[7][96] 	= partial_clause_prev[7][96] & ~x[37];
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & ~x[39];
			partial_clause[7][99] 	= partial_clause_prev[7][99] & ~x[39];
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & x[16];
			partial_clause[8][1] 	= partial_clause_prev[8][1] & x[17];
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & x[16];
			partial_clause[8][4] 	= partial_clause_prev[8][4] & x[17] & ~x[56];
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & x[18];
			partial_clause[8][7] 	= partial_clause_prev[8][7] & x[16];
			partial_clause[8][8] 	= partial_clause_prev[8][8] & x[16];
			partial_clause[8][9] 	= partial_clause_prev[8][9] & x[15];
			partial_clause[8][10] 	= partial_clause_prev[8][10] & x[15] & ~x[36];
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & x[17];
			partial_clause[8][14] 	= partial_clause_prev[8][14] & x[17] & ~x[32];
			partial_clause[8][15] 	= partial_clause_prev[8][15] & ~x[3] & x[16];
			partial_clause[8][16] 	= partial_clause_prev[8][16] & x[17] & ~x[31] & ~x[32];
			partial_clause[8][17] 	= partial_clause_prev[8][17] & x[17];
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & x[16] & ~x[27];
			partial_clause[8][20] 	= partial_clause_prev[8][20] & x[16] & x[18];
			partial_clause[8][21] 	= partial_clause_prev[8][21] & x[16];
			partial_clause[8][22] 	= partial_clause_prev[8][22] & x[16];
			partial_clause[8][23] 	= partial_clause_prev[8][23] & x[16];
			partial_clause[8][24] 	= partial_clause_prev[8][24] & x[17];
			partial_clause[8][25] 	= partial_clause_prev[8][25] & x[16];
			partial_clause[8][26] 	= partial_clause_prev[8][26] & x[16];
			partial_clause[8][27] 	= partial_clause_prev[8][27] & x[16];
			partial_clause[8][28] 	= partial_clause_prev[8][28] & ~x[5] & x[17] & ~x[33];
			partial_clause[8][29] 	= partial_clause_prev[8][29] & x[16];
			partial_clause[8][30] 	= partial_clause_prev[8][30] & x[16];
			partial_clause[8][31] 	= partial_clause_prev[8][31] & x[17] & ~x[58];
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & ~x[36];
			partial_clause[8][35] 	= partial_clause_prev[8][35] & x[17] & ~x[58];
			partial_clause[8][36] 	= partial_clause_prev[8][36] & x[16];
			partial_clause[8][37] 	= partial_clause_prev[8][37] & x[16] & x[17];
			partial_clause[8][38] 	= partial_clause_prev[8][38] & x[18] & ~x[57];
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & x[17];
			partial_clause[8][41] 	= partial_clause_prev[8][41] & x[15] & ~x[33];
			partial_clause[8][42] 	= partial_clause_prev[8][42] & x[15];
			partial_clause[8][43] 	= partial_clause_prev[8][43] & x[16];
			partial_clause[8][44] 	= partial_clause_prev[8][44] & ~x[5] & x[17];
			partial_clause[8][45] 	= partial_clause_prev[8][45] & ~x[26];
			partial_clause[8][46] 	= partial_clause_prev[8][46] & ~x[27];
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & x[17];
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & ~x[59];
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & ~x[21] & ~x[46];
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & ~x[14];
			partial_clause[8][56] 	= partial_clause_prev[8][56] & ~x[1];
			partial_clause[8][57] 	= partial_clause_prev[8][57] & ~x[3];
			partial_clause[8][58] 	= partial_clause_prev[8][58] & ~x[5] & ~x[24];
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & ~x[24];
			partial_clause[8][61] 	= partial_clause_prev[8][61] & ~x[18] & ~x[45];
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & ~x[12] & ~x[13] & ~x[19];
			partial_clause[8][64] 	= partial_clause_prev[8][64] & ~x[23] & ~x[32];
			partial_clause[8][65] 	= partial_clause_prev[8][65] & ~x[4] & ~x[15] & ~x[20];
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & ~x[30];
			partial_clause[8][69] 	= partial_clause_prev[8][69] & ~x[13] & ~x[20] & ~x[27] & ~x[41];
			partial_clause[8][70] 	= partial_clause_prev[8][70] & ~x[32];
			partial_clause[8][71] 	= partial_clause_prev[8][71] & ~x[33];
			partial_clause[8][72] 	= partial_clause_prev[8][72] & ~x[12] & ~x[18] & ~x[46];
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & ~x[29];
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & ~x[58];
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & ~x[36];
			partial_clause[8][81] 	= partial_clause_prev[8][81] & ~x[4] & ~x[16] & ~x[20] & ~x[43];
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & ~x[39] & ~x[54];
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & ~x[13] & ~x[14] & ~x[20] & ~x[48];
			partial_clause[8][86] 	= partial_clause_prev[8][86] & ~x[0] & ~x[4];
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & ~x[53];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & ~x[16] & ~x[17] & ~x[18];
			partial_clause[8][92] 	= partial_clause_prev[8][92] & ~x[17] & ~x[45];
			partial_clause[8][93] 	= partial_clause_prev[8][93] & ~x[55] & ~x[59];
			partial_clause[8][94] 	= partial_clause_prev[8][94] & ~x[2];
			partial_clause[8][95] 	= partial_clause_prev[8][95] & ~x[14] & ~x[31] & ~x[40];
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & ~x[12];
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & ~x[14];
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & ~x[12] & ~x[40];
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & ~x[11];
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & ~x[10];
			partial_clause[9][36] 	= partial_clause_prev[9][36] & ~x[10];
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & ~x[13];
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & ~x[26] & ~x[49];
			partial_clause[9][51] 	= partial_clause_prev[9][51] & ~x[29];
			partial_clause[9][52] 	= partial_clause_prev[9][52] & ~x[6];
			partial_clause[9][53] 	= partial_clause_prev[9][53] & 1'b1;
			partial_clause[9][54] 	= partial_clause_prev[9][54] & ~x[52];
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & ~x[50] & ~x[51];
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & ~x[49] & ~x[51];
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & ~x[1];
			partial_clause[9][61] 	= partial_clause_prev[9][61] & ~x[34] & ~x[52];
			partial_clause[9][62] 	= partial_clause_prev[9][62] & ~x[50];
			partial_clause[9][63] 	= partial_clause_prev[9][63] & ~x[40] & ~x[51];
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & ~x[47] & ~x[50];
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & ~x[51] & ~x[58];
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & ~x[2] & ~x[51] & ~x[52];
			partial_clause[9][70] 	= partial_clause_prev[9][70] & ~x[55];
			partial_clause[9][71] 	= partial_clause_prev[9][71] & ~x[49];
			partial_clause[9][72] 	= partial_clause_prev[9][72] & ~x[29];
			partial_clause[9][73] 	= partial_clause_prev[9][73] & ~x[52];
			partial_clause[9][74] 	= partial_clause_prev[9][74] & ~x[37] & ~x[56];
			partial_clause[9][75] 	= partial_clause_prev[9][75] & ~x[51] & ~x[52];
			partial_clause[9][76] 	= partial_clause_prev[9][76] & ~x[46] & ~x[50] & ~x[52];
			partial_clause[9][77] 	= partial_clause_prev[9][77] & ~x[49] & ~x[50];
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & ~x[51];
			partial_clause[9][81] 	= partial_clause_prev[9][81] & ~x[39] & ~x[44] & ~x[50] & ~x[52];
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & 1'b1;
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & ~x[26] & ~x[49];
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & ~x[49] & ~x[51];
			partial_clause[9][90] 	= partial_clause_prev[9][90] & ~x[61];
			partial_clause[9][91] 	= partial_clause_prev[9][91] & ~x[53];
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & ~x[24] & ~x[26] & ~x[50];
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & ~x[48] & ~x[50];
			partial_clause[9][97] 	= partial_clause_prev[9][97] & ~x[2] & ~x[24] & ~x[25] & ~x[50];
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & ~x[52];
		end
	end
endmodule


module HCB_11 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & ~x[38];
			partial_clause[0][1] 	= partial_clause_prev[0][1] & ~x[31];
			partial_clause[0][2] 	= partial_clause_prev[0][2] & ~x[6] & ~x[7];
			partial_clause[0][3] 	= partial_clause_prev[0][3] & ~x[57];
			partial_clause[0][4] 	= partial_clause_prev[0][4] & ~x[11];
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & ~x[38];
			partial_clause[0][7] 	= partial_clause_prev[0][7] & ~x[8] & ~x[53];
			partial_clause[0][8] 	= partial_clause_prev[0][8] & ~x[10];
			partial_clause[0][9] 	= partial_clause_prev[0][9] & ~x[14] & ~x[20];
			partial_clause[0][10] 	= partial_clause_prev[0][10] & ~x[13] & ~x[36] & ~x[40];
			partial_clause[0][11] 	= partial_clause_prev[0][11] & ~x[9] & ~x[11] & ~x[57];
			partial_clause[0][12] 	= partial_clause_prev[0][12] & ~x[6] & ~x[7];
			partial_clause[0][13] 	= partial_clause_prev[0][13] & ~x[6] & ~x[11] & ~x[35];
			partial_clause[0][14] 	= partial_clause_prev[0][14] & ~x[8];
			partial_clause[0][15] 	= partial_clause_prev[0][15] & ~x[35];
			partial_clause[0][16] 	= partial_clause_prev[0][16] & ~x[5] & ~x[15] & ~x[37];
			partial_clause[0][17] 	= partial_clause_prev[0][17] & ~x[12];
			partial_clause[0][18] 	= partial_clause_prev[0][18] & ~x[7] & ~x[39];
			partial_clause[0][19] 	= partial_clause_prev[0][19] & 1'b1;
			partial_clause[0][20] 	= partial_clause_prev[0][20] & ~x[51];
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & ~x[36];
			partial_clause[0][23] 	= partial_clause_prev[0][23] & ~x[9];
			partial_clause[0][24] 	= partial_clause_prev[0][24] & ~x[60];
			partial_clause[0][25] 	= partial_clause_prev[0][25] & ~x[10] & ~x[35] & ~x[62];
			partial_clause[0][26] 	= partial_clause_prev[0][26] & ~x[6] & ~x[19] & ~x[37];
			partial_clause[0][27] 	= partial_clause_prev[0][27] & ~x[8] & ~x[11] & ~x[39];
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & ~x[4] & ~x[37];
			partial_clause[0][30] 	= partial_clause_prev[0][30] & ~x[8];
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & ~x[12] & ~x[38];
			partial_clause[0][33] 	= partial_clause_prev[0][33] & ~x[7] & ~x[18];
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & ~x[7] & ~x[39];
			partial_clause[0][36] 	= partial_clause_prev[0][36] & ~x[38] & ~x[58];
			partial_clause[0][37] 	= partial_clause_prev[0][37] & ~x[38] & ~x[40];
			partial_clause[0][38] 	= partial_clause_prev[0][38] & ~x[13];
			partial_clause[0][39] 	= partial_clause_prev[0][39] & ~x[17];
			partial_clause[0][40] 	= partial_clause_prev[0][40] & ~x[10];
			partial_clause[0][41] 	= partial_clause_prev[0][41] & ~x[13];
			partial_clause[0][42] 	= partial_clause_prev[0][42] & 1'b1;
			partial_clause[0][43] 	= partial_clause_prev[0][43] & 1'b1;
			partial_clause[0][44] 	= partial_clause_prev[0][44] & ~x[10];
			partial_clause[0][45] 	= partial_clause_prev[0][45] & ~x[4] & ~x[10] & ~x[54];
			partial_clause[0][46] 	= partial_clause_prev[0][46] & ~x[7];
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & ~x[10];
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & 1'b1;
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & ~x[24];
			partial_clause[0][53] 	= partial_clause_prev[0][53] & 1'b1;
			partial_clause[0][54] 	= partial_clause_prev[0][54] & ~x[60];
			partial_clause[0][55] 	= partial_clause_prev[0][55] & ~x[52];
			partial_clause[0][56] 	= partial_clause_prev[0][56] & ~x[19];
			partial_clause[0][57] 	= partial_clause_prev[0][57] & ~x[48] & ~x[49];
			partial_clause[0][58] 	= partial_clause_prev[0][58] & ~x[23] & ~x[51];
			partial_clause[0][59] 	= partial_clause_prev[0][59] & ~x[54];
			partial_clause[0][60] 	= partial_clause_prev[0][60] & 1'b1;
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & 1'b1;
			partial_clause[0][64] 	= partial_clause_prev[0][64] & ~x[21] & ~x[22] & ~x[29];
			partial_clause[0][65] 	= partial_clause_prev[0][65] & ~x[20] & ~x[55];
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & ~x[48];
			partial_clause[0][68] 	= partial_clause_prev[0][68] & 1'b1;
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & ~x[23] & ~x[44];
			partial_clause[0][71] 	= partial_clause_prev[0][71] & ~x[42];
			partial_clause[0][72] 	= partial_clause_prev[0][72] & ~x[18] & ~x[19] & ~x[45];
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & ~x[1];
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & ~x[48];
			partial_clause[0][78] 	= partial_clause_prev[0][78] & 1'b1;
			partial_clause[0][79] 	= partial_clause_prev[0][79] & ~x[17];
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & ~x[51];
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & ~x[23] & ~x[43];
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & ~x[45];
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & ~x[17];
			partial_clause[0][91] 	= partial_clause_prev[0][91] & ~x[31];
			partial_clause[0][92] 	= partial_clause_prev[0][92] & 1'b1;
			partial_clause[0][93] 	= partial_clause_prev[0][93] & ~x[48];
			partial_clause[0][94] 	= partial_clause_prev[0][94] & ~x[56];
			partial_clause[0][95] 	= partial_clause_prev[0][95] & 1'b1;
			partial_clause[0][96] 	= partial_clause_prev[0][96] & ~x[20] & ~x[25];
			partial_clause[0][97] 	= partial_clause_prev[0][97] & ~x[0] & ~x[22] & ~x[52];
			partial_clause[0][98] 	= partial_clause_prev[0][98] & 1'b1;
			partial_clause[0][99] 	= partial_clause_prev[0][99] & ~x[47];
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & ~x[6];
			partial_clause[1][10] 	= partial_clause_prev[1][10] & ~x[54];
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & ~x[25];
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & ~x[6];
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & ~x[57];
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & ~x[6];
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & ~x[8];
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & ~x[49];
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & ~x[0] & ~x[22];
			partial_clause[1][52] 	= partial_clause_prev[1][52] & ~x[25];
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & ~x[59];
			partial_clause[1][55] 	= partial_clause_prev[1][55] & ~x[54];
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & ~x[2];
			partial_clause[1][58] 	= partial_clause_prev[1][58] & 1'b1;
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & ~x[1] & ~x[16] & ~x[62];
			partial_clause[1][61] 	= partial_clause_prev[1][61] & ~x[24] & ~x[47];
			partial_clause[1][62] 	= partial_clause_prev[1][62] & ~x[1] & ~x[47] & ~x[53];
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & ~x[30] & ~x[51];
			partial_clause[1][65] 	= partial_clause_prev[1][65] & ~x[40] & ~x[48];
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & ~x[18] & ~x[54];
			partial_clause[1][69] 	= partial_clause_prev[1][69] & ~x[24] & ~x[47] & ~x[61];
			partial_clause[1][70] 	= partial_clause_prev[1][70] & ~x[21] & ~x[24] & ~x[50];
			partial_clause[1][71] 	= partial_clause_prev[1][71] & 1'b1;
			partial_clause[1][72] 	= partial_clause_prev[1][72] & 1'b1;
			partial_clause[1][73] 	= partial_clause_prev[1][73] & ~x[50];
			partial_clause[1][74] 	= partial_clause_prev[1][74] & ~x[63];
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & 1'b1;
			partial_clause[1][77] 	= partial_clause_prev[1][77] & ~x[28];
			partial_clause[1][78] 	= partial_clause_prev[1][78] & ~x[51];
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & ~x[48];
			partial_clause[1][81] 	= partial_clause_prev[1][81] & ~x[41];
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & ~x[46];
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & ~x[29] & ~x[51];
			partial_clause[1][86] 	= partial_clause_prev[1][86] & ~x[2];
			partial_clause[1][87] 	= partial_clause_prev[1][87] & ~x[30];
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & ~x[60];
			partial_clause[1][90] 	= partial_clause_prev[1][90] & 1'b1;
			partial_clause[1][91] 	= partial_clause_prev[1][91] & ~x[31];
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & ~x[45];
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & ~x[26];
			partial_clause[1][97] 	= partial_clause_prev[1][97] & ~x[20];
			partial_clause[1][98] 	= partial_clause_prev[1][98] & ~x[20] & ~x[42] & ~x[43];
			partial_clause[1][99] 	= partial_clause_prev[1][99] & ~x[54];
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & ~x[44];
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & ~x[3];
			partial_clause[2][4] 	= partial_clause_prev[2][4] & ~x[26] & ~x[40];
			partial_clause[2][5] 	= partial_clause_prev[2][5] & 1'b1;
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & ~x[2];
			partial_clause[2][8] 	= partial_clause_prev[2][8] & ~x[8];
			partial_clause[2][9] 	= partial_clause_prev[2][9] & ~x[21] & ~x[28];
			partial_clause[2][10] 	= partial_clause_prev[2][10] & ~x[9] & ~x[22];
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & ~x[11] & ~x[14] & ~x[60];
			partial_clause[2][16] 	= partial_clause_prev[2][16] & ~x[11];
			partial_clause[2][17] 	= partial_clause_prev[2][17] & ~x[6] & ~x[10];
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & ~x[47];
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & ~x[38] & ~x[48];
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & ~x[40];
			partial_clause[2][26] 	= partial_clause_prev[2][26] & ~x[23];
			partial_clause[2][27] 	= partial_clause_prev[2][27] & ~x[13];
			partial_clause[2][28] 	= partial_clause_prev[2][28] & ~x[62];
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & ~x[8];
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & 1'b1;
			partial_clause[2][33] 	= partial_clause_prev[2][33] & 1'b1;
			partial_clause[2][34] 	= partial_clause_prev[2][34] & ~x[7];
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & ~x[11] & ~x[36];
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & ~x[31];
			partial_clause[2][41] 	= partial_clause_prev[2][41] & ~x[0];
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & ~x[5];
			partial_clause[2][44] 	= partial_clause_prev[2][44] & ~x[47];
			partial_clause[2][45] 	= partial_clause_prev[2][45] & ~x[5] & ~x[11];
			partial_clause[2][46] 	= partial_clause_prev[2][46] & ~x[38] & ~x[48];
			partial_clause[2][47] 	= partial_clause_prev[2][47] & ~x[31];
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & 1'b1;
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & ~x[56] & ~x[59];
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & ~x[19];
			partial_clause[2][64] 	= partial_clause_prev[2][64] & ~x[49] & ~x[61];
			partial_clause[2][65] 	= partial_clause_prev[2][65] & ~x[51];
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & ~x[60];
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & ~x[18];
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & ~x[53];
			partial_clause[2][80] 	= partial_clause_prev[2][80] & 1'b1;
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & ~x[52];
			partial_clause[2][85] 	= partial_clause_prev[2][85] & 1'b1;
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & ~x[51] & ~x[63];
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & ~x[0];
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & ~x[48];
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & ~x[52];
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & ~x[48];
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & ~x[37];
			partial_clause[3][1] 	= partial_clause_prev[3][1] & ~x[10];
			partial_clause[3][2] 	= partial_clause_prev[3][2] & ~x[12] & ~x[52];
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & ~x[32];
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & ~x[36];
			partial_clause[3][9] 	= partial_clause_prev[3][9] & 1'b1;
			partial_clause[3][10] 	= partial_clause_prev[3][10] & ~x[40];
			partial_clause[3][11] 	= partial_clause_prev[3][11] & 1'b1;
			partial_clause[3][12] 	= partial_clause_prev[3][12] & ~x[39];
			partial_clause[3][13] 	= partial_clause_prev[3][13] & ~x[26];
			partial_clause[3][14] 	= partial_clause_prev[3][14] & 1'b1;
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & ~x[51];
			partial_clause[3][19] 	= partial_clause_prev[3][19] & 1'b1;
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & ~x[12] & ~x[35];
			partial_clause[3][24] 	= partial_clause_prev[3][24] & ~x[37];
			partial_clause[3][25] 	= partial_clause_prev[3][25] & ~x[13];
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & ~x[18];
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & 1'b1;
			partial_clause[3][30] 	= partial_clause_prev[3][30] & ~x[32];
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & ~x[21];
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & ~x[28] & ~x[48];
			partial_clause[3][40] 	= partial_clause_prev[3][40] & ~x[38];
			partial_clause[3][41] 	= partial_clause_prev[3][41] & ~x[50];
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & ~x[38];
			partial_clause[3][47] 	= partial_clause_prev[3][47] & ~x[35] & ~x[49];
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & 1'b1;
			partial_clause[3][51] 	= partial_clause_prev[3][51] & ~x[3] & ~x[48];
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & ~x[27];
			partial_clause[3][55] 	= partial_clause_prev[3][55] & ~x[8];
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & ~x[29] & ~x[46] & ~x[54];
			partial_clause[3][60] 	= partial_clause_prev[3][60] & 1'b1;
			partial_clause[3][61] 	= partial_clause_prev[3][61] & ~x[46];
			partial_clause[3][62] 	= partial_clause_prev[3][62] & 1'b1;
			partial_clause[3][63] 	= partial_clause_prev[3][63] & ~x[46];
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[22];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & ~x[24];
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & ~x[20];
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & ~x[51];
			partial_clause[3][72] 	= partial_clause_prev[3][72] & ~x[50];
			partial_clause[3][73] 	= partial_clause_prev[3][73] & ~x[38];
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & ~x[22];
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & ~x[21];
			partial_clause[3][79] 	= partial_clause_prev[3][79] & ~x[30];
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & ~x[54];
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & ~x[20];
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & ~x[3];
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & ~x[23];
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & ~x[44];
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & ~x[16];
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & ~x[38] & ~x[46];
			partial_clause[4][1] 	= partial_clause_prev[4][1] & ~x[35];
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & ~x[2] & ~x[34];
			partial_clause[4][4] 	= partial_clause_prev[4][4] & ~x[38];
			partial_clause[4][5] 	= partial_clause_prev[4][5] & 1'b1;
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & ~x[61];
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & ~x[4];
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & ~x[34];
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & ~x[7];
			partial_clause[4][15] 	= partial_clause_prev[4][15] & ~x[35];
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & ~x[36];
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & ~x[37];
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & ~x[44];
			partial_clause[4][25] 	= partial_clause_prev[4][25] & ~x[39] & ~x[41];
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & ~x[25];
			partial_clause[4][32] 	= partial_clause_prev[4][32] & ~x[3];
			partial_clause[4][33] 	= partial_clause_prev[4][33] & 1'b1;
			partial_clause[4][34] 	= partial_clause_prev[4][34] & ~x[35] & ~x[37] & ~x[41];
			partial_clause[4][35] 	= partial_clause_prev[4][35] & ~x[5];
			partial_clause[4][36] 	= partial_clause_prev[4][36] & ~x[54];
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & ~x[37] & ~x[39];
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & ~x[8] & ~x[35] & ~x[40];
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & 1'b1;
			partial_clause[4][50] 	= partial_clause_prev[4][50] & 1'b1;
			partial_clause[4][51] 	= partial_clause_prev[4][51] & 1'b1;
			partial_clause[4][52] 	= partial_clause_prev[4][52] & ~x[27];
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & ~x[55] & ~x[61];
			partial_clause[4][55] 	= partial_clause_prev[4][55] & ~x[28] & ~x[50];
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & ~x[28] & ~x[29];
			partial_clause[4][58] 	= partial_clause_prev[4][58] & ~x[22];
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & 1'b1;
			partial_clause[4][61] 	= partial_clause_prev[4][61] & ~x[39];
			partial_clause[4][62] 	= partial_clause_prev[4][62] & ~x[25] & ~x[26];
			partial_clause[4][63] 	= partial_clause_prev[4][63] & ~x[58];
			partial_clause[4][64] 	= partial_clause_prev[4][64] & 1'b1;
			partial_clause[4][65] 	= partial_clause_prev[4][65] & ~x[24];
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & ~x[21] & ~x[44] & ~x[52];
			partial_clause[4][68] 	= partial_clause_prev[4][68] & 1'b1;
			partial_clause[4][69] 	= partial_clause_prev[4][69] & ~x[52];
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & ~x[51] & ~x[60];
			partial_clause[4][72] 	= partial_clause_prev[4][72] & ~x[17];
			partial_clause[4][73] 	= partial_clause_prev[4][73] & 1'b1;
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & ~x[26];
			partial_clause[4][77] 	= partial_clause_prev[4][77] & ~x[57];
			partial_clause[4][78] 	= partial_clause_prev[4][78] & ~x[18] & ~x[26];
			partial_clause[4][79] 	= partial_clause_prev[4][79] & 1'b1;
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & ~x[1] & ~x[26];
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & ~x[50];
			partial_clause[4][86] 	= partial_clause_prev[4][86] & ~x[21];
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & ~x[48];
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & ~x[56];
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & ~x[23] & ~x[25];
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & ~x[31] & ~x[45];
			partial_clause[4][97] 	= partial_clause_prev[4][97] & 1'b1;
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & ~x[34];
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & ~x[50];
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & ~x[22];
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & ~x[0];
			partial_clause[5][11] 	= partial_clause_prev[5][11] & ~x[17];
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & ~x[37];
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & ~x[31] & ~x[33];
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & ~x[16];
			partial_clause[5][23] 	= partial_clause_prev[5][23] & ~x[26] & ~x[36];
			partial_clause[5][24] 	= partial_clause_prev[5][24] & ~x[51] & ~x[57];
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & ~x[48];
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & 1'b1;
			partial_clause[5][43] 	= partial_clause_prev[5][43] & ~x[27];
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & ~x[35] & ~x[38];
			partial_clause[5][48] 	= partial_clause_prev[5][48] & ~x[31];
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & ~x[43];
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & 1'b1;
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & ~x[55];
			partial_clause[5][67] 	= partial_clause_prev[5][67] & ~x[21];
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & ~x[23];
			partial_clause[5][71] 	= partial_clause_prev[5][71] & ~x[44];
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & 1'b1;
			partial_clause[5][75] 	= partial_clause_prev[5][75] & ~x[28];
			partial_clause[5][76] 	= partial_clause_prev[5][76] & ~x[40];
			partial_clause[5][77] 	= partial_clause_prev[5][77] & ~x[47];
			partial_clause[5][78] 	= partial_clause_prev[5][78] & 1'b1;
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & ~x[0];
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & ~x[45];
			partial_clause[5][90] 	= partial_clause_prev[5][90] & 1'b1;
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & ~x[58];
			partial_clause[5][96] 	= partial_clause_prev[5][96] & ~x[15];
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & ~x[27] & ~x[49] & ~x[61];
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & 1'b1;
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & 1'b1;
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & ~x[38];
			partial_clause[6][7] 	= partial_clause_prev[6][7] & ~x[7] & ~x[30];
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & ~x[29];
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & ~x[61];
			partial_clause[6][12] 	= partial_clause_prev[6][12] & ~x[48];
			partial_clause[6][13] 	= partial_clause_prev[6][13] & ~x[44];
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & ~x[3];
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & ~x[13] & ~x[37];
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & ~x[10];
			partial_clause[6][22] 	= partial_clause_prev[6][22] & ~x[7];
			partial_clause[6][23] 	= partial_clause_prev[6][23] & ~x[8];
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & ~x[40];
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & ~x[38] & ~x[56];
			partial_clause[6][36] 	= partial_clause_prev[6][36] & ~x[23];
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & ~x[6];
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & ~x[57];
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & ~x[26];
			partial_clause[6][56] 	= partial_clause_prev[6][56] & ~x[2];
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & ~x[44];
			partial_clause[6][60] 	= partial_clause_prev[6][60] & ~x[56];
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & ~x[20];
			partial_clause[6][64] 	= partial_clause_prev[6][64] & ~x[20] & ~x[21];
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & ~x[19];
			partial_clause[6][70] 	= partial_clause_prev[6][70] & ~x[56];
			partial_clause[6][71] 	= partial_clause_prev[6][71] & ~x[62];
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & 1'b1;
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & ~x[49];
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & ~x[20];
			partial_clause[6][83] 	= partial_clause_prev[6][83] & ~x[27];
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & ~x[44] & ~x[63];
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & ~x[21];
			partial_clause[6][91] 	= partial_clause_prev[6][91] & 1'b1;
			partial_clause[6][92] 	= partial_clause_prev[6][92] & ~x[21] & ~x[51];
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & ~x[23];
			partial_clause[6][96] 	= partial_clause_prev[6][96] & 1'b1;
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & ~x[27];
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & ~x[46];
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & ~x[56];
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & ~x[57];
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & ~x[45];
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & ~x[5];
			partial_clause[7][51] 	= partial_clause_prev[7][51] & ~x[3] & ~x[5] & ~x[6] & ~x[8] & ~x[10] & ~x[39] & ~x[41];
			partial_clause[7][52] 	= partial_clause_prev[7][52] & ~x[5] & ~x[7] & ~x[10] & ~x[12] & ~x[36];
			partial_clause[7][53] 	= partial_clause_prev[7][53] & ~x[23] & ~x[32];
			partial_clause[7][54] 	= partial_clause_prev[7][54] & ~x[4] & ~x[5] & ~x[9] & ~x[11];
			partial_clause[7][55] 	= partial_clause_prev[7][55] & ~x[5] & ~x[7] & ~x[8] & ~x[11];
			partial_clause[7][56] 	= partial_clause_prev[7][56] & ~x[10] & ~x[33];
			partial_clause[7][57] 	= partial_clause_prev[7][57] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[13];
			partial_clause[7][58] 	= partial_clause_prev[7][58] & ~x[5] & ~x[7] & ~x[8] & ~x[10] & ~x[13];
			partial_clause[7][59] 	= partial_clause_prev[7][59] & ~x[6] & ~x[9] & ~x[10] & ~x[11] & ~x[12];
			partial_clause[7][60] 	= partial_clause_prev[7][60] & ~x[3] & ~x[5] & ~x[7] & ~x[11] & ~x[13];
			partial_clause[7][61] 	= partial_clause_prev[7][61] & ~x[7] & ~x[11] & ~x[13] & ~x[32] & ~x[33] & ~x[41];
			partial_clause[7][62] 	= partial_clause_prev[7][62] & ~x[8] & ~x[10] & ~x[11] & ~x[40];
			partial_clause[7][63] 	= partial_clause_prev[7][63] & ~x[58] & ~x[61];
			partial_clause[7][64] 	= partial_clause_prev[7][64] & ~x[3] & ~x[6] & ~x[7] & ~x[8] & ~x[11] & ~x[41];
			partial_clause[7][65] 	= partial_clause_prev[7][65] & ~x[4] & ~x[7] & ~x[8] & ~x[10] & ~x[40];
			partial_clause[7][66] 	= partial_clause_prev[7][66] & ~x[5] & ~x[8] & ~x[11] & ~x[12] & ~x[33];
			partial_clause[7][67] 	= partial_clause_prev[7][67] & ~x[1] & ~x[5] & ~x[7] & ~x[9] & ~x[10] & ~x[11] & ~x[42];
			partial_clause[7][68] 	= partial_clause_prev[7][68] & ~x[15] & ~x[37];
			partial_clause[7][69] 	= partial_clause_prev[7][69] & ~x[6] & ~x[8] & ~x[12] & ~x[39];
			partial_clause[7][70] 	= partial_clause_prev[7][70] & ~x[5] & ~x[7] & ~x[9] & ~x[11] & ~x[13];
			partial_clause[7][71] 	= partial_clause_prev[7][71] & ~x[15] & ~x[25] & ~x[38];
			partial_clause[7][72] 	= partial_clause_prev[7][72] & ~x[4] & ~x[5] & ~x[6] & ~x[8] & ~x[10] & ~x[12] & ~x[18];
			partial_clause[7][73] 	= partial_clause_prev[7][73] & ~x[6] & ~x[9] & ~x[10];
			partial_clause[7][74] 	= partial_clause_prev[7][74] & ~x[3] & ~x[6] & ~x[7] & ~x[10] & ~x[13];
			partial_clause[7][75] 	= partial_clause_prev[7][75] & ~x[6] & ~x[9] & ~x[39];
			partial_clause[7][76] 	= partial_clause_prev[7][76] & ~x[2] & ~x[4] & ~x[5] & ~x[7] & ~x[9] & ~x[10] & ~x[11];
			partial_clause[7][77] 	= partial_clause_prev[7][77] & ~x[2] & ~x[4] & ~x[7] & ~x[9];
			partial_clause[7][78] 	= partial_clause_prev[7][78] & ~x[6] & ~x[7] & ~x[9] & ~x[11] & ~x[12] & ~x[49];
			partial_clause[7][79] 	= partial_clause_prev[7][79] & ~x[19];
			partial_clause[7][80] 	= partial_clause_prev[7][80] & ~x[5] & ~x[6] & ~x[11] & ~x[35] & ~x[56];
			partial_clause[7][81] 	= partial_clause_prev[7][81] & ~x[5] & ~x[7] & ~x[9] & ~x[10] & ~x[12] & ~x[13] & ~x[49];
			partial_clause[7][82] 	= partial_clause_prev[7][82] & ~x[38] & ~x[47];
			partial_clause[7][83] 	= partial_clause_prev[7][83] & ~x[4] & ~x[8] & ~x[11] & ~x[36] & ~x[58];
			partial_clause[7][84] 	= partial_clause_prev[7][84] & ~x[3] & ~x[5] & ~x[7] & ~x[10] & ~x[11] & ~x[13] & ~x[33];
			partial_clause[7][85] 	= partial_clause_prev[7][85] & ~x[5] & ~x[7] & ~x[9] & ~x[10] & ~x[13] & ~x[63];
			partial_clause[7][86] 	= partial_clause_prev[7][86] & ~x[33] & ~x[34] & ~x[37];
			partial_clause[7][87] 	= partial_clause_prev[7][87] & ~x[4] & ~x[7] & ~x[8] & ~x[10] & ~x[11] & ~x[12];
			partial_clause[7][88] 	= partial_clause_prev[7][88] & ~x[7] & ~x[9] & ~x[11] & ~x[12] & ~x[41];
			partial_clause[7][89] 	= partial_clause_prev[7][89] & ~x[7] & ~x[28];
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & ~x[6];
			partial_clause[7][92] 	= partial_clause_prev[7][92] & ~x[4] & ~x[5] & ~x[6] & ~x[8] & ~x[9] & ~x[34];
			partial_clause[7][93] 	= partial_clause_prev[7][93] & ~x[3] & ~x[5] & ~x[6] & ~x[8] & ~x[10];
			partial_clause[7][94] 	= partial_clause_prev[7][94] & ~x[27] & ~x[39] & ~x[45] & ~x[48] & ~x[49];
			partial_clause[7][95] 	= partial_clause_prev[7][95] & ~x[4] & ~x[7] & ~x[9] & ~x[15];
			partial_clause[7][96] 	= partial_clause_prev[7][96] & ~x[5] & ~x[7] & ~x[9] & ~x[13] & ~x[41];
			partial_clause[7][97] 	= partial_clause_prev[7][97] & ~x[4] & ~x[5] & ~x[6] & ~x[8] & ~x[10] & ~x[12] & ~x[36];
			partial_clause[7][98] 	= partial_clause_prev[7][98] & ~x[4] & ~x[7] & ~x[9] & ~x[39] & ~x[57];
			partial_clause[7][99] 	= partial_clause_prev[7][99] & ~x[2] & ~x[5] & ~x[6] & ~x[7] & ~x[9] & ~x[10] & ~x[12];
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & ~x[36];
			partial_clause[8][1] 	= partial_clause_prev[8][1] & 1'b1;
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & ~x[2] & ~x[32];
			partial_clause[8][4] 	= partial_clause_prev[8][4] & ~x[22];
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & ~x[28];
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & ~x[39];
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & ~x[51];
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & ~x[25];
			partial_clause[8][18] 	= partial_clause_prev[8][18] & ~x[36];
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & 1'b1;
			partial_clause[8][22] 	= partial_clause_prev[8][22] & ~x[19] & ~x[26];
			partial_clause[8][23] 	= partial_clause_prev[8][23] & ~x[30];
			partial_clause[8][24] 	= partial_clause_prev[8][24] & ~x[20] & ~x[54];
			partial_clause[8][25] 	= partial_clause_prev[8][25] & ~x[53];
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & ~x[8];
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & ~x[3];
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & ~x[28];
			partial_clause[8][32] 	= partial_clause_prev[8][32] & 1'b1;
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & ~x[19];
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & ~x[0] & ~x[26];
			partial_clause[8][38] 	= partial_clause_prev[8][38] & ~x[34];
			partial_clause[8][39] 	= partial_clause_prev[8][39] & ~x[3];
			partial_clause[8][40] 	= partial_clause_prev[8][40] & ~x[23];
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & ~x[40];
			partial_clause[8][43] 	= partial_clause_prev[8][43] & ~x[45];
			partial_clause[8][44] 	= partial_clause_prev[8][44] & 1'b1;
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & 1'b1;
			partial_clause[8][47] 	= partial_clause_prev[8][47] & ~x[25] & ~x[38] & ~x[49] & ~x[54];
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & ~x[35] & ~x[42];
			partial_clause[8][50] 	= partial_clause_prev[8][50] & 1'b1;
			partial_clause[8][51] 	= partial_clause_prev[8][51] & 1'b1;
			partial_clause[8][52] 	= partial_clause_prev[8][52] & ~x[6];
			partial_clause[8][53] 	= partial_clause_prev[8][53] & 1'b1;
			partial_clause[8][54] 	= partial_clause_prev[8][54] & 1'b1;
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & ~x[22];
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & ~x[24];
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & 1'b1;
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & ~x[51];
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & ~x[28];
			partial_clause[8][68] 	= partial_clause_prev[8][68] & ~x[22];
			partial_clause[8][69] 	= partial_clause_prev[8][69] & ~x[51];
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & ~x[22] & ~x[56];
			partial_clause[8][72] 	= partial_clause_prev[8][72] & ~x[61];
			partial_clause[8][73] 	= partial_clause_prev[8][73] & ~x[50];
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & ~x[55];
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & ~x[55];
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & ~x[22] & ~x[45] & ~x[55];
			partial_clause[8][84] 	= partial_clause_prev[8][84] & 1'b1;
			partial_clause[8][85] 	= partial_clause_prev[8][85] & ~x[62];
			partial_clause[8][86] 	= partial_clause_prev[8][86] & ~x[18] & ~x[59];
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & ~x[46];
			partial_clause[8][89] 	= partial_clause_prev[8][89] & ~x[48];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & 1'b1;
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & ~x[27];
			partial_clause[8][94] 	= partial_clause_prev[8][94] & 1'b1;
			partial_clause[8][95] 	= partial_clause_prev[8][95] & 1'b1;
			partial_clause[8][96] 	= partial_clause_prev[8][96] & 1'b1;
			partial_clause[8][97] 	= partial_clause_prev[8][97] & ~x[1];
			partial_clause[8][98] 	= partial_clause_prev[8][98] & ~x[27] & ~x[43];
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & ~x[47];
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & ~x[21];
			partial_clause[9][8] 	= partial_clause_prev[9][8] & ~x[59];
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & 1'b1;
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & 1'b1;
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & 1'b1;
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & ~x[45];
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & 1'b1;
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & ~x[58];
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & ~x[3] & ~x[5] & ~x[7] & ~x[8] & ~x[10] & ~x[11] & ~x[42];
			partial_clause[9][51] 	= partial_clause_prev[9][51] & ~x[4] & ~x[8] & ~x[9];
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & ~x[4] & ~x[6] & ~x[7] & ~x[9] & ~x[36];
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & ~x[4] & ~x[5] & ~x[43];
			partial_clause[9][56] 	= partial_clause_prev[9][56] & ~x[38] & ~x[40];
			partial_clause[9][57] 	= partial_clause_prev[9][57] & ~x[4] & ~x[16];
			partial_clause[9][58] 	= partial_clause_prev[9][58] & ~x[4] & ~x[6] & ~x[10] & ~x[11] & ~x[12];
			partial_clause[9][59] 	= partial_clause_prev[9][59] & ~x[17] & ~x[44] & ~x[60];
			partial_clause[9][60] 	= partial_clause_prev[9][60] & ~x[4] & ~x[6] & ~x[55];
			partial_clause[9][61] 	= partial_clause_prev[9][61] & ~x[9] & ~x[10] & ~x[11] & ~x[13] & ~x[15];
			partial_clause[9][62] 	= partial_clause_prev[9][62] & ~x[5] & ~x[7] & ~x[9] & ~x[11] & ~x[13] & ~x[15];
			partial_clause[9][63] 	= partial_clause_prev[9][63] & ~x[0] & ~x[6] & ~x[8] & ~x[11] & ~x[13] & ~x[34];
			partial_clause[9][64] 	= partial_clause_prev[9][64] & ~x[3] & ~x[4] & ~x[15] & ~x[16];
			partial_clause[9][65] 	= partial_clause_prev[9][65] & ~x[5] & ~x[6] & ~x[10] & ~x[14] & ~x[15] & ~x[17] & ~x[39];
			partial_clause[9][66] 	= partial_clause_prev[9][66] & ~x[3];
			partial_clause[9][67] 	= partial_clause_prev[9][67] & ~x[10] & ~x[11] & ~x[12] & ~x[15];
			partial_clause[9][68] 	= partial_clause_prev[9][68] & ~x[13] & ~x[19] & ~x[38];
			partial_clause[9][69] 	= partial_clause_prev[9][69] & ~x[14];
			partial_clause[9][70] 	= partial_clause_prev[9][70] & ~x[5] & ~x[49] & ~x[61];
			partial_clause[9][71] 	= partial_clause_prev[9][71] & ~x[4] & ~x[5] & ~x[7] & ~x[9] & ~x[10] & ~x[11] & ~x[14] & ~x[16];
			partial_clause[9][72] 	= partial_clause_prev[9][72] & ~x[3] & ~x[6] & ~x[7] & ~x[16];
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & ~x[57];
			partial_clause[9][75] 	= partial_clause_prev[9][75] & ~x[4] & ~x[6] & ~x[13] & ~x[14];
			partial_clause[9][76] 	= partial_clause_prev[9][76] & ~x[4] & ~x[9] & ~x[10] & ~x[12];
			partial_clause[9][77] 	= partial_clause_prev[9][77] & ~x[6] & ~x[8] & ~x[9] & ~x[51];
			partial_clause[9][78] 	= partial_clause_prev[9][78] & ~x[57];
			partial_clause[9][79] 	= partial_clause_prev[9][79] & ~x[8] & ~x[10] & ~x[11] & ~x[13] & ~x[15] & ~x[36] & ~x[48];
			partial_clause[9][80] 	= partial_clause_prev[9][80] & ~x[3] & ~x[6] & ~x[7] & ~x[9] & ~x[10] & ~x[12] & ~x[14] & ~x[62];
			partial_clause[9][81] 	= partial_clause_prev[9][81] & ~x[7] & ~x[10] & ~x[11] & ~x[12] & ~x[13];
			partial_clause[9][82] 	= partial_clause_prev[9][82] & ~x[1] & ~x[5] & ~x[7] & ~x[14];
			partial_clause[9][83] 	= partial_clause_prev[9][83] & ~x[8] & ~x[10];
			partial_clause[9][84] 	= partial_clause_prev[9][84] & ~x[4] & ~x[5] & ~x[7] & ~x[11] & ~x[13] & ~x[17] & ~x[34];
			partial_clause[9][85] 	= partial_clause_prev[9][85] & ~x[2] & ~x[6] & ~x[8] & ~x[9] & ~x[11];
			partial_clause[9][86] 	= partial_clause_prev[9][86] & ~x[4] & ~x[6];
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & ~x[3] & ~x[5] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[16];
			partial_clause[9][90] 	= partial_clause_prev[9][90] & ~x[7] & ~x[51];
			partial_clause[9][91] 	= partial_clause_prev[9][91] & ~x[4];
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & ~x[11];
			partial_clause[9][94] 	= partial_clause_prev[9][94] & ~x[4] & ~x[6] & ~x[9] & ~x[10] & ~x[12];
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & ~x[5] & ~x[7] & ~x[9] & ~x[10] & ~x[12] & ~x[42];
			partial_clause[9][97] 	= partial_clause_prev[9][97] & ~x[5] & ~x[6] & ~x[9] & ~x[11] & ~x[12];
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & ~x[7] & ~x[10] & ~x[13] & ~x[58];
		end
	end
endmodule


module HCB_12 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [99:0] partial_clause_prev [10];
	output	logic[99:0] partial_clause [10];
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			// Class 0
			partial_clause[0][0] 	= partial_clause_prev[0][0] & 1'b1;
			partial_clause[0][1] 	= partial_clause_prev[0][1] & 1'b1;
			partial_clause[0][2] 	= partial_clause_prev[0][2] & 1'b1;
			partial_clause[0][3] 	= partial_clause_prev[0][3] & 1'b1;
			partial_clause[0][4] 	= partial_clause_prev[0][4] & 1'b1;
			partial_clause[0][5] 	= partial_clause_prev[0][5] & 1'b1;
			partial_clause[0][6] 	= partial_clause_prev[0][6] & 1'b1;
			partial_clause[0][7] 	= partial_clause_prev[0][7] & 1'b1;
			partial_clause[0][8] 	= partial_clause_prev[0][8] & 1'b1;
			partial_clause[0][9] 	= partial_clause_prev[0][9] & 1'b1;
			partial_clause[0][10] 	= partial_clause_prev[0][10] & 1'b1;
			partial_clause[0][11] 	= partial_clause_prev[0][11] & 1'b1;
			partial_clause[0][12] 	= partial_clause_prev[0][12] & 1'b1;
			partial_clause[0][13] 	= partial_clause_prev[0][13] & 1'b1;
			partial_clause[0][14] 	= partial_clause_prev[0][14] & 1'b1;
			partial_clause[0][15] 	= partial_clause_prev[0][15] & 1'b1;
			partial_clause[0][16] 	= partial_clause_prev[0][16] & 1'b1;
			partial_clause[0][17] 	= partial_clause_prev[0][17] & 1'b1;
			partial_clause[0][18] 	= partial_clause_prev[0][18] & 1'b1;
			partial_clause[0][19] 	= partial_clause_prev[0][19] & ~x[4];
			partial_clause[0][20] 	= partial_clause_prev[0][20] & 1'b1;
			partial_clause[0][21] 	= partial_clause_prev[0][21] & 1'b1;
			partial_clause[0][22] 	= partial_clause_prev[0][22] & 1'b1;
			partial_clause[0][23] 	= partial_clause_prev[0][23] & 1'b1;
			partial_clause[0][24] 	= partial_clause_prev[0][24] & 1'b1;
			partial_clause[0][25] 	= partial_clause_prev[0][25] & 1'b1;
			partial_clause[0][26] 	= partial_clause_prev[0][26] & 1'b1;
			partial_clause[0][27] 	= partial_clause_prev[0][27] & 1'b1;
			partial_clause[0][28] 	= partial_clause_prev[0][28] & 1'b1;
			partial_clause[0][29] 	= partial_clause_prev[0][29] & ~x[12];
			partial_clause[0][30] 	= partial_clause_prev[0][30] & ~x[4];
			partial_clause[0][31] 	= partial_clause_prev[0][31] & 1'b1;
			partial_clause[0][32] 	= partial_clause_prev[0][32] & 1'b1;
			partial_clause[0][33] 	= partial_clause_prev[0][33] & 1'b1;
			partial_clause[0][34] 	= partial_clause_prev[0][34] & 1'b1;
			partial_clause[0][35] 	= partial_clause_prev[0][35] & 1'b1;
			partial_clause[0][36] 	= partial_clause_prev[0][36] & 1'b1;
			partial_clause[0][37] 	= partial_clause_prev[0][37] & 1'b1;
			partial_clause[0][38] 	= partial_clause_prev[0][38] & 1'b1;
			partial_clause[0][39] 	= partial_clause_prev[0][39] & ~x[3];
			partial_clause[0][40] 	= partial_clause_prev[0][40] & 1'b1;
			partial_clause[0][41] 	= partial_clause_prev[0][41] & 1'b1;
			partial_clause[0][42] 	= partial_clause_prev[0][42] & ~x[5] & ~x[12];
			partial_clause[0][43] 	= partial_clause_prev[0][43] & ~x[1];
			partial_clause[0][44] 	= partial_clause_prev[0][44] & 1'b1;
			partial_clause[0][45] 	= partial_clause_prev[0][45] & 1'b1;
			partial_clause[0][46] 	= partial_clause_prev[0][46] & 1'b1;
			partial_clause[0][47] 	= partial_clause_prev[0][47] & 1'b1;
			partial_clause[0][48] 	= partial_clause_prev[0][48] & 1'b1;
			partial_clause[0][49] 	= partial_clause_prev[0][49] & 1'b1;
			partial_clause[0][50] 	= partial_clause_prev[0][50] & ~x[15];
			partial_clause[0][51] 	= partial_clause_prev[0][51] & 1'b1;
			partial_clause[0][52] 	= partial_clause_prev[0][52] & 1'b1;
			partial_clause[0][53] 	= partial_clause_prev[0][53] & ~x[13];
			partial_clause[0][54] 	= partial_clause_prev[0][54] & 1'b1;
			partial_clause[0][55] 	= partial_clause_prev[0][55] & 1'b1;
			partial_clause[0][56] 	= partial_clause_prev[0][56] & ~x[1];
			partial_clause[0][57] 	= partial_clause_prev[0][57] & 1'b1;
			partial_clause[0][58] 	= partial_clause_prev[0][58] & 1'b1;
			partial_clause[0][59] 	= partial_clause_prev[0][59] & 1'b1;
			partial_clause[0][60] 	= partial_clause_prev[0][60] & ~x[4] & ~x[5];
			partial_clause[0][61] 	= partial_clause_prev[0][61] & 1'b1;
			partial_clause[0][62] 	= partial_clause_prev[0][62] & 1'b1;
			partial_clause[0][63] 	= partial_clause_prev[0][63] & ~x[4];
			partial_clause[0][64] 	= partial_clause_prev[0][64] & 1'b1;
			partial_clause[0][65] 	= partial_clause_prev[0][65] & 1'b1;
			partial_clause[0][66] 	= partial_clause_prev[0][66] & 1'b1;
			partial_clause[0][67] 	= partial_clause_prev[0][67] & 1'b1;
			partial_clause[0][68] 	= partial_clause_prev[0][68] & ~x[3] & ~x[12];
			partial_clause[0][69] 	= partial_clause_prev[0][69] & 1'b1;
			partial_clause[0][70] 	= partial_clause_prev[0][70] & 1'b1;
			partial_clause[0][71] 	= partial_clause_prev[0][71] & 1'b1;
			partial_clause[0][72] 	= partial_clause_prev[0][72] & ~x[4];
			partial_clause[0][73] 	= partial_clause_prev[0][73] & 1'b1;
			partial_clause[0][74] 	= partial_clause_prev[0][74] & 1'b1;
			partial_clause[0][75] 	= partial_clause_prev[0][75] & 1'b1;
			partial_clause[0][76] 	= partial_clause_prev[0][76] & 1'b1;
			partial_clause[0][77] 	= partial_clause_prev[0][77] & 1'b1;
			partial_clause[0][78] 	= partial_clause_prev[0][78] & ~x[5];
			partial_clause[0][79] 	= partial_clause_prev[0][79] & 1'b1;
			partial_clause[0][80] 	= partial_clause_prev[0][80] & 1'b1;
			partial_clause[0][81] 	= partial_clause_prev[0][81] & 1'b1;
			partial_clause[0][82] 	= partial_clause_prev[0][82] & 1'b1;
			partial_clause[0][83] 	= partial_clause_prev[0][83] & 1'b1;
			partial_clause[0][84] 	= partial_clause_prev[0][84] & 1'b1;
			partial_clause[0][85] 	= partial_clause_prev[0][85] & 1'b1;
			partial_clause[0][86] 	= partial_clause_prev[0][86] & 1'b1;
			partial_clause[0][87] 	= partial_clause_prev[0][87] & 1'b1;
			partial_clause[0][88] 	= partial_clause_prev[0][88] & ~x[8] & ~x[12];
			partial_clause[0][89] 	= partial_clause_prev[0][89] & 1'b1;
			partial_clause[0][90] 	= partial_clause_prev[0][90] & ~x[4];
			partial_clause[0][91] 	= partial_clause_prev[0][91] & ~x[7];
			partial_clause[0][92] 	= partial_clause_prev[0][92] & ~x[7];
			partial_clause[0][93] 	= partial_clause_prev[0][93] & 1'b1;
			partial_clause[0][94] 	= partial_clause_prev[0][94] & ~x[13];
			partial_clause[0][95] 	= partial_clause_prev[0][95] & ~x[0];
			partial_clause[0][96] 	= partial_clause_prev[0][96] & ~x[15];
			partial_clause[0][97] 	= partial_clause_prev[0][97] & 1'b1;
			partial_clause[0][98] 	= partial_clause_prev[0][98] & ~x[1];
			partial_clause[0][99] 	= partial_clause_prev[0][99] & 1'b1;
			// Class 1
			partial_clause[1][0] 	= partial_clause_prev[1][0] & 1'b1;
			partial_clause[1][1] 	= partial_clause_prev[1][1] & 1'b1;
			partial_clause[1][2] 	= partial_clause_prev[1][2] & 1'b1;
			partial_clause[1][3] 	= partial_clause_prev[1][3] & 1'b1;
			partial_clause[1][4] 	= partial_clause_prev[1][4] & 1'b1;
			partial_clause[1][5] 	= partial_clause_prev[1][5] & 1'b1;
			partial_clause[1][6] 	= partial_clause_prev[1][6] & 1'b1;
			partial_clause[1][7] 	= partial_clause_prev[1][7] & 1'b1;
			partial_clause[1][8] 	= partial_clause_prev[1][8] & 1'b1;
			partial_clause[1][9] 	= partial_clause_prev[1][9] & 1'b1;
			partial_clause[1][10] 	= partial_clause_prev[1][10] & 1'b1;
			partial_clause[1][11] 	= partial_clause_prev[1][11] & 1'b1;
			partial_clause[1][12] 	= partial_clause_prev[1][12] & 1'b1;
			partial_clause[1][13] 	= partial_clause_prev[1][13] & 1'b1;
			partial_clause[1][14] 	= partial_clause_prev[1][14] & 1'b1;
			partial_clause[1][15] 	= partial_clause_prev[1][15] & 1'b1;
			partial_clause[1][16] 	= partial_clause_prev[1][16] & 1'b1;
			partial_clause[1][17] 	= partial_clause_prev[1][17] & 1'b1;
			partial_clause[1][18] 	= partial_clause_prev[1][18] & 1'b1;
			partial_clause[1][19] 	= partial_clause_prev[1][19] & 1'b1;
			partial_clause[1][20] 	= partial_clause_prev[1][20] & 1'b1;
			partial_clause[1][21] 	= partial_clause_prev[1][21] & 1'b1;
			partial_clause[1][22] 	= partial_clause_prev[1][22] & 1'b1;
			partial_clause[1][23] 	= partial_clause_prev[1][23] & 1'b1;
			partial_clause[1][24] 	= partial_clause_prev[1][24] & 1'b1;
			partial_clause[1][25] 	= partial_clause_prev[1][25] & 1'b1;
			partial_clause[1][26] 	= partial_clause_prev[1][26] & 1'b1;
			partial_clause[1][27] 	= partial_clause_prev[1][27] & 1'b1;
			partial_clause[1][28] 	= partial_clause_prev[1][28] & 1'b1;
			partial_clause[1][29] 	= partial_clause_prev[1][29] & 1'b1;
			partial_clause[1][30] 	= partial_clause_prev[1][30] & 1'b1;
			partial_clause[1][31] 	= partial_clause_prev[1][31] & 1'b1;
			partial_clause[1][32] 	= partial_clause_prev[1][32] & 1'b1;
			partial_clause[1][33] 	= partial_clause_prev[1][33] & 1'b1;
			partial_clause[1][34] 	= partial_clause_prev[1][34] & 1'b1;
			partial_clause[1][35] 	= partial_clause_prev[1][35] & 1'b1;
			partial_clause[1][36] 	= partial_clause_prev[1][36] & 1'b1;
			partial_clause[1][37] 	= partial_clause_prev[1][37] & 1'b1;
			partial_clause[1][38] 	= partial_clause_prev[1][38] & 1'b1;
			partial_clause[1][39] 	= partial_clause_prev[1][39] & 1'b1;
			partial_clause[1][40] 	= partial_clause_prev[1][40] & 1'b1;
			partial_clause[1][41] 	= partial_clause_prev[1][41] & 1'b1;
			partial_clause[1][42] 	= partial_clause_prev[1][42] & 1'b1;
			partial_clause[1][43] 	= partial_clause_prev[1][43] & 1'b1;
			partial_clause[1][44] 	= partial_clause_prev[1][44] & 1'b1;
			partial_clause[1][45] 	= partial_clause_prev[1][45] & 1'b1;
			partial_clause[1][46] 	= partial_clause_prev[1][46] & 1'b1;
			partial_clause[1][47] 	= partial_clause_prev[1][47] & 1'b1;
			partial_clause[1][48] 	= partial_clause_prev[1][48] & 1'b1;
			partial_clause[1][49] 	= partial_clause_prev[1][49] & 1'b1;
			partial_clause[1][50] 	= partial_clause_prev[1][50] & 1'b1;
			partial_clause[1][51] 	= partial_clause_prev[1][51] & 1'b1;
			partial_clause[1][52] 	= partial_clause_prev[1][52] & 1'b1;
			partial_clause[1][53] 	= partial_clause_prev[1][53] & 1'b1;
			partial_clause[1][54] 	= partial_clause_prev[1][54] & 1'b1;
			partial_clause[1][55] 	= partial_clause_prev[1][55] & 1'b1;
			partial_clause[1][56] 	= partial_clause_prev[1][56] & 1'b1;
			partial_clause[1][57] 	= partial_clause_prev[1][57] & 1'b1;
			partial_clause[1][58] 	= partial_clause_prev[1][58] & 1'b1;
			partial_clause[1][59] 	= partial_clause_prev[1][59] & 1'b1;
			partial_clause[1][60] 	= partial_clause_prev[1][60] & 1'b1;
			partial_clause[1][61] 	= partial_clause_prev[1][61] & ~x[10];
			partial_clause[1][62] 	= partial_clause_prev[1][62] & ~x[14];
			partial_clause[1][63] 	= partial_clause_prev[1][63] & 1'b1;
			partial_clause[1][64] 	= partial_clause_prev[1][64] & ~x[15];
			partial_clause[1][65] 	= partial_clause_prev[1][65] & 1'b1;
			partial_clause[1][66] 	= partial_clause_prev[1][66] & 1'b1;
			partial_clause[1][67] 	= partial_clause_prev[1][67] & 1'b1;
			partial_clause[1][68] 	= partial_clause_prev[1][68] & ~x[15];
			partial_clause[1][69] 	= partial_clause_prev[1][69] & 1'b1;
			partial_clause[1][70] 	= partial_clause_prev[1][70] & ~x[6] & ~x[15];
			partial_clause[1][71] 	= partial_clause_prev[1][71] & ~x[11] & ~x[15];
			partial_clause[1][72] 	= partial_clause_prev[1][72] & ~x[12];
			partial_clause[1][73] 	= partial_clause_prev[1][73] & ~x[12];
			partial_clause[1][74] 	= partial_clause_prev[1][74] & 1'b1;
			partial_clause[1][75] 	= partial_clause_prev[1][75] & 1'b1;
			partial_clause[1][76] 	= partial_clause_prev[1][76] & ~x[6];
			partial_clause[1][77] 	= partial_clause_prev[1][77] & 1'b1;
			partial_clause[1][78] 	= partial_clause_prev[1][78] & 1'b1;
			partial_clause[1][79] 	= partial_clause_prev[1][79] & 1'b1;
			partial_clause[1][80] 	= partial_clause_prev[1][80] & 1'b1;
			partial_clause[1][81] 	= partial_clause_prev[1][81] & ~x[13];
			partial_clause[1][82] 	= partial_clause_prev[1][82] & 1'b1;
			partial_clause[1][83] 	= partial_clause_prev[1][83] & 1'b1;
			partial_clause[1][84] 	= partial_clause_prev[1][84] & 1'b1;
			partial_clause[1][85] 	= partial_clause_prev[1][85] & 1'b1;
			partial_clause[1][86] 	= partial_clause_prev[1][86] & 1'b1;
			partial_clause[1][87] 	= partial_clause_prev[1][87] & 1'b1;
			partial_clause[1][88] 	= partial_clause_prev[1][88] & 1'b1;
			partial_clause[1][89] 	= partial_clause_prev[1][89] & 1'b1;
			partial_clause[1][90] 	= partial_clause_prev[1][90] & ~x[6];
			partial_clause[1][91] 	= partial_clause_prev[1][91] & 1'b1;
			partial_clause[1][92] 	= partial_clause_prev[1][92] & 1'b1;
			partial_clause[1][93] 	= partial_clause_prev[1][93] & ~x[10];
			partial_clause[1][94] 	= partial_clause_prev[1][94] & 1'b1;
			partial_clause[1][95] 	= partial_clause_prev[1][95] & 1'b1;
			partial_clause[1][96] 	= partial_clause_prev[1][96] & 1'b1;
			partial_clause[1][97] 	= partial_clause_prev[1][97] & ~x[8];
			partial_clause[1][98] 	= partial_clause_prev[1][98] & 1'b1;
			partial_clause[1][99] 	= partial_clause_prev[1][99] & 1'b1;
			// Class 2
			partial_clause[2][0] 	= partial_clause_prev[2][0] & 1'b1;
			partial_clause[2][1] 	= partial_clause_prev[2][1] & 1'b1;
			partial_clause[2][2] 	= partial_clause_prev[2][2] & 1'b1;
			partial_clause[2][3] 	= partial_clause_prev[2][3] & 1'b1;
			partial_clause[2][4] 	= partial_clause_prev[2][4] & 1'b1;
			partial_clause[2][5] 	= partial_clause_prev[2][5] & ~x[1] & ~x[11];
			partial_clause[2][6] 	= partial_clause_prev[2][6] & 1'b1;
			partial_clause[2][7] 	= partial_clause_prev[2][7] & ~x[15];
			partial_clause[2][8] 	= partial_clause_prev[2][8] & 1'b1;
			partial_clause[2][9] 	= partial_clause_prev[2][9] & 1'b1;
			partial_clause[2][10] 	= partial_clause_prev[2][10] & 1'b1;
			partial_clause[2][11] 	= partial_clause_prev[2][11] & 1'b1;
			partial_clause[2][12] 	= partial_clause_prev[2][12] & 1'b1;
			partial_clause[2][13] 	= partial_clause_prev[2][13] & 1'b1;
			partial_clause[2][14] 	= partial_clause_prev[2][14] & 1'b1;
			partial_clause[2][15] 	= partial_clause_prev[2][15] & 1'b1;
			partial_clause[2][16] 	= partial_clause_prev[2][16] & 1'b1;
			partial_clause[2][17] 	= partial_clause_prev[2][17] & 1'b1;
			partial_clause[2][18] 	= partial_clause_prev[2][18] & 1'b1;
			partial_clause[2][19] 	= partial_clause_prev[2][19] & 1'b1;
			partial_clause[2][20] 	= partial_clause_prev[2][20] & 1'b1;
			partial_clause[2][21] 	= partial_clause_prev[2][21] & 1'b1;
			partial_clause[2][22] 	= partial_clause_prev[2][22] & 1'b1;
			partial_clause[2][23] 	= partial_clause_prev[2][23] & 1'b1;
			partial_clause[2][24] 	= partial_clause_prev[2][24] & 1'b1;
			partial_clause[2][25] 	= partial_clause_prev[2][25] & 1'b1;
			partial_clause[2][26] 	= partial_clause_prev[2][26] & 1'b1;
			partial_clause[2][27] 	= partial_clause_prev[2][27] & 1'b1;
			partial_clause[2][28] 	= partial_clause_prev[2][28] & 1'b1;
			partial_clause[2][29] 	= partial_clause_prev[2][29] & 1'b1;
			partial_clause[2][30] 	= partial_clause_prev[2][30] & 1'b1;
			partial_clause[2][31] 	= partial_clause_prev[2][31] & 1'b1;
			partial_clause[2][32] 	= partial_clause_prev[2][32] & ~x[9];
			partial_clause[2][33] 	= partial_clause_prev[2][33] & ~x[15];
			partial_clause[2][34] 	= partial_clause_prev[2][34] & 1'b1;
			partial_clause[2][35] 	= partial_clause_prev[2][35] & 1'b1;
			partial_clause[2][36] 	= partial_clause_prev[2][36] & 1'b1;
			partial_clause[2][37] 	= partial_clause_prev[2][37] & 1'b1;
			partial_clause[2][38] 	= partial_clause_prev[2][38] & 1'b1;
			partial_clause[2][39] 	= partial_clause_prev[2][39] & 1'b1;
			partial_clause[2][40] 	= partial_clause_prev[2][40] & 1'b1;
			partial_clause[2][41] 	= partial_clause_prev[2][41] & 1'b1;
			partial_clause[2][42] 	= partial_clause_prev[2][42] & 1'b1;
			partial_clause[2][43] 	= partial_clause_prev[2][43] & ~x[5];
			partial_clause[2][44] 	= partial_clause_prev[2][44] & 1'b1;
			partial_clause[2][45] 	= partial_clause_prev[2][45] & 1'b1;
			partial_clause[2][46] 	= partial_clause_prev[2][46] & 1'b1;
			partial_clause[2][47] 	= partial_clause_prev[2][47] & 1'b1;
			partial_clause[2][48] 	= partial_clause_prev[2][48] & 1'b1;
			partial_clause[2][49] 	= partial_clause_prev[2][49] & ~x[12] & ~x[14];
			partial_clause[2][50] 	= partial_clause_prev[2][50] & 1'b1;
			partial_clause[2][51] 	= partial_clause_prev[2][51] & 1'b1;
			partial_clause[2][52] 	= partial_clause_prev[2][52] & 1'b1;
			partial_clause[2][53] 	= partial_clause_prev[2][53] & 1'b1;
			partial_clause[2][54] 	= partial_clause_prev[2][54] & 1'b1;
			partial_clause[2][55] 	= partial_clause_prev[2][55] & 1'b1;
			partial_clause[2][56] 	= partial_clause_prev[2][56] & 1'b1;
			partial_clause[2][57] 	= partial_clause_prev[2][57] & 1'b1;
			partial_clause[2][58] 	= partial_clause_prev[2][58] & 1'b1;
			partial_clause[2][59] 	= partial_clause_prev[2][59] & 1'b1;
			partial_clause[2][60] 	= partial_clause_prev[2][60] & 1'b1;
			partial_clause[2][61] 	= partial_clause_prev[2][61] & 1'b1;
			partial_clause[2][62] 	= partial_clause_prev[2][62] & 1'b1;
			partial_clause[2][63] 	= partial_clause_prev[2][63] & 1'b1;
			partial_clause[2][64] 	= partial_clause_prev[2][64] & 1'b1;
			partial_clause[2][65] 	= partial_clause_prev[2][65] & 1'b1;
			partial_clause[2][66] 	= partial_clause_prev[2][66] & 1'b1;
			partial_clause[2][67] 	= partial_clause_prev[2][67] & 1'b1;
			partial_clause[2][68] 	= partial_clause_prev[2][68] & 1'b1;
			partial_clause[2][69] 	= partial_clause_prev[2][69] & 1'b1;
			partial_clause[2][70] 	= partial_clause_prev[2][70] & 1'b1;
			partial_clause[2][71] 	= partial_clause_prev[2][71] & 1'b1;
			partial_clause[2][72] 	= partial_clause_prev[2][72] & 1'b1;
			partial_clause[2][73] 	= partial_clause_prev[2][73] & 1'b1;
			partial_clause[2][74] 	= partial_clause_prev[2][74] & 1'b1;
			partial_clause[2][75] 	= partial_clause_prev[2][75] & 1'b1;
			partial_clause[2][76] 	= partial_clause_prev[2][76] & 1'b1;
			partial_clause[2][77] 	= partial_clause_prev[2][77] & 1'b1;
			partial_clause[2][78] 	= partial_clause_prev[2][78] & 1'b1;
			partial_clause[2][79] 	= partial_clause_prev[2][79] & 1'b1;
			partial_clause[2][80] 	= partial_clause_prev[2][80] & ~x[11];
			partial_clause[2][81] 	= partial_clause_prev[2][81] & 1'b1;
			partial_clause[2][82] 	= partial_clause_prev[2][82] & 1'b1;
			partial_clause[2][83] 	= partial_clause_prev[2][83] & 1'b1;
			partial_clause[2][84] 	= partial_clause_prev[2][84] & 1'b1;
			partial_clause[2][85] 	= partial_clause_prev[2][85] & ~x[13];
			partial_clause[2][86] 	= partial_clause_prev[2][86] & 1'b1;
			partial_clause[2][87] 	= partial_clause_prev[2][87] & 1'b1;
			partial_clause[2][88] 	= partial_clause_prev[2][88] & 1'b1;
			partial_clause[2][89] 	= partial_clause_prev[2][89] & 1'b1;
			partial_clause[2][90] 	= partial_clause_prev[2][90] & 1'b1;
			partial_clause[2][91] 	= partial_clause_prev[2][91] & 1'b1;
			partial_clause[2][92] 	= partial_clause_prev[2][92] & 1'b1;
			partial_clause[2][93] 	= partial_clause_prev[2][93] & 1'b1;
			partial_clause[2][94] 	= partial_clause_prev[2][94] & 1'b1;
			partial_clause[2][95] 	= partial_clause_prev[2][95] & 1'b1;
			partial_clause[2][96] 	= partial_clause_prev[2][96] & 1'b1;
			partial_clause[2][97] 	= partial_clause_prev[2][97] & 1'b1;
			partial_clause[2][98] 	= partial_clause_prev[2][98] & 1'b1;
			partial_clause[2][99] 	= partial_clause_prev[2][99] & 1'b1;
			// Class 3
			partial_clause[3][0] 	= partial_clause_prev[3][0] & 1'b1;
			partial_clause[3][1] 	= partial_clause_prev[3][1] & 1'b1;
			partial_clause[3][2] 	= partial_clause_prev[3][2] & 1'b1;
			partial_clause[3][3] 	= partial_clause_prev[3][3] & 1'b1;
			partial_clause[3][4] 	= partial_clause_prev[3][4] & 1'b1;
			partial_clause[3][5] 	= partial_clause_prev[3][5] & 1'b1;
			partial_clause[3][6] 	= partial_clause_prev[3][6] & 1'b1;
			partial_clause[3][7] 	= partial_clause_prev[3][7] & 1'b1;
			partial_clause[3][8] 	= partial_clause_prev[3][8] & 1'b1;
			partial_clause[3][9] 	= partial_clause_prev[3][9] & ~x[9];
			partial_clause[3][10] 	= partial_clause_prev[3][10] & 1'b1;
			partial_clause[3][11] 	= partial_clause_prev[3][11] & ~x[0];
			partial_clause[3][12] 	= partial_clause_prev[3][12] & 1'b1;
			partial_clause[3][13] 	= partial_clause_prev[3][13] & 1'b1;
			partial_clause[3][14] 	= partial_clause_prev[3][14] & ~x[12];
			partial_clause[3][15] 	= partial_clause_prev[3][15] & 1'b1;
			partial_clause[3][16] 	= partial_clause_prev[3][16] & 1'b1;
			partial_clause[3][17] 	= partial_clause_prev[3][17] & 1'b1;
			partial_clause[3][18] 	= partial_clause_prev[3][18] & 1'b1;
			partial_clause[3][19] 	= partial_clause_prev[3][19] & ~x[15];
			partial_clause[3][20] 	= partial_clause_prev[3][20] & 1'b1;
			partial_clause[3][21] 	= partial_clause_prev[3][21] & 1'b1;
			partial_clause[3][22] 	= partial_clause_prev[3][22] & 1'b1;
			partial_clause[3][23] 	= partial_clause_prev[3][23] & ~x[8];
			partial_clause[3][24] 	= partial_clause_prev[3][24] & 1'b1;
			partial_clause[3][25] 	= partial_clause_prev[3][25] & 1'b1;
			partial_clause[3][26] 	= partial_clause_prev[3][26] & 1'b1;
			partial_clause[3][27] 	= partial_clause_prev[3][27] & 1'b1;
			partial_clause[3][28] 	= partial_clause_prev[3][28] & 1'b1;
			partial_clause[3][29] 	= partial_clause_prev[3][29] & ~x[6];
			partial_clause[3][30] 	= partial_clause_prev[3][30] & 1'b1;
			partial_clause[3][31] 	= partial_clause_prev[3][31] & 1'b1;
			partial_clause[3][32] 	= partial_clause_prev[3][32] & 1'b1;
			partial_clause[3][33] 	= partial_clause_prev[3][33] & 1'b1;
			partial_clause[3][34] 	= partial_clause_prev[3][34] & 1'b1;
			partial_clause[3][35] 	= partial_clause_prev[3][35] & 1'b1;
			partial_clause[3][36] 	= partial_clause_prev[3][36] & 1'b1;
			partial_clause[3][37] 	= partial_clause_prev[3][37] & 1'b1;
			partial_clause[3][38] 	= partial_clause_prev[3][38] & 1'b1;
			partial_clause[3][39] 	= partial_clause_prev[3][39] & 1'b1;
			partial_clause[3][40] 	= partial_clause_prev[3][40] & 1'b1;
			partial_clause[3][41] 	= partial_clause_prev[3][41] & 1'b1;
			partial_clause[3][42] 	= partial_clause_prev[3][42] & 1'b1;
			partial_clause[3][43] 	= partial_clause_prev[3][43] & 1'b1;
			partial_clause[3][44] 	= partial_clause_prev[3][44] & 1'b1;
			partial_clause[3][45] 	= partial_clause_prev[3][45] & 1'b1;
			partial_clause[3][46] 	= partial_clause_prev[3][46] & 1'b1;
			partial_clause[3][47] 	= partial_clause_prev[3][47] & 1'b1;
			partial_clause[3][48] 	= partial_clause_prev[3][48] & 1'b1;
			partial_clause[3][49] 	= partial_clause_prev[3][49] & 1'b1;
			partial_clause[3][50] 	= partial_clause_prev[3][50] & ~x[7] & ~x[13];
			partial_clause[3][51] 	= partial_clause_prev[3][51] & 1'b1;
			partial_clause[3][52] 	= partial_clause_prev[3][52] & 1'b1;
			partial_clause[3][53] 	= partial_clause_prev[3][53] & 1'b1;
			partial_clause[3][54] 	= partial_clause_prev[3][54] & 1'b1;
			partial_clause[3][55] 	= partial_clause_prev[3][55] & ~x[9];
			partial_clause[3][56] 	= partial_clause_prev[3][56] & 1'b1;
			partial_clause[3][57] 	= partial_clause_prev[3][57] & 1'b1;
			partial_clause[3][58] 	= partial_clause_prev[3][58] & 1'b1;
			partial_clause[3][59] 	= partial_clause_prev[3][59] & 1'b1;
			partial_clause[3][60] 	= partial_clause_prev[3][60] & ~x[0];
			partial_clause[3][61] 	= partial_clause_prev[3][61] & 1'b1;
			partial_clause[3][62] 	= partial_clause_prev[3][62] & ~x[5];
			partial_clause[3][63] 	= partial_clause_prev[3][63] & ~x[10];
			partial_clause[3][64] 	= partial_clause_prev[3][64] & 1'b1;
			partial_clause[3][65] 	= partial_clause_prev[3][65] & ~x[12];
			partial_clause[3][66] 	= partial_clause_prev[3][66] & 1'b1;
			partial_clause[3][67] 	= partial_clause_prev[3][67] & 1'b1;
			partial_clause[3][68] 	= partial_clause_prev[3][68] & 1'b1;
			partial_clause[3][69] 	= partial_clause_prev[3][69] & 1'b1;
			partial_clause[3][70] 	= partial_clause_prev[3][70] & 1'b1;
			partial_clause[3][71] 	= partial_clause_prev[3][71] & 1'b1;
			partial_clause[3][72] 	= partial_clause_prev[3][72] & 1'b1;
			partial_clause[3][73] 	= partial_clause_prev[3][73] & 1'b1;
			partial_clause[3][74] 	= partial_clause_prev[3][74] & 1'b1;
			partial_clause[3][75] 	= partial_clause_prev[3][75] & 1'b1;
			partial_clause[3][76] 	= partial_clause_prev[3][76] & 1'b1;
			partial_clause[3][77] 	= partial_clause_prev[3][77] & 1'b1;
			partial_clause[3][78] 	= partial_clause_prev[3][78] & 1'b1;
			partial_clause[3][79] 	= partial_clause_prev[3][79] & 1'b1;
			partial_clause[3][80] 	= partial_clause_prev[3][80] & 1'b1;
			partial_clause[3][81] 	= partial_clause_prev[3][81] & 1'b1;
			partial_clause[3][82] 	= partial_clause_prev[3][82] & 1'b1;
			partial_clause[3][83] 	= partial_clause_prev[3][83] & 1'b1;
			partial_clause[3][84] 	= partial_clause_prev[3][84] & 1'b1;
			partial_clause[3][85] 	= partial_clause_prev[3][85] & 1'b1;
			partial_clause[3][86] 	= partial_clause_prev[3][86] & 1'b1;
			partial_clause[3][87] 	= partial_clause_prev[3][87] & 1'b1;
			partial_clause[3][88] 	= partial_clause_prev[3][88] & 1'b1;
			partial_clause[3][89] 	= partial_clause_prev[3][89] & 1'b1;
			partial_clause[3][90] 	= partial_clause_prev[3][90] & 1'b1;
			partial_clause[3][91] 	= partial_clause_prev[3][91] & 1'b1;
			partial_clause[3][92] 	= partial_clause_prev[3][92] & 1'b1;
			partial_clause[3][93] 	= partial_clause_prev[3][93] & 1'b1;
			partial_clause[3][94] 	= partial_clause_prev[3][94] & 1'b1;
			partial_clause[3][95] 	= partial_clause_prev[3][95] & 1'b1;
			partial_clause[3][96] 	= partial_clause_prev[3][96] & 1'b1;
			partial_clause[3][97] 	= partial_clause_prev[3][97] & 1'b1;
			partial_clause[3][98] 	= partial_clause_prev[3][98] & 1'b1;
			partial_clause[3][99] 	= partial_clause_prev[3][99] & 1'b1;
			// Class 4
			partial_clause[4][0] 	= partial_clause_prev[4][0] & 1'b1;
			partial_clause[4][1] 	= partial_clause_prev[4][1] & 1'b1;
			partial_clause[4][2] 	= partial_clause_prev[4][2] & 1'b1;
			partial_clause[4][3] 	= partial_clause_prev[4][3] & 1'b1;
			partial_clause[4][4] 	= partial_clause_prev[4][4] & 1'b1;
			partial_clause[4][5] 	= partial_clause_prev[4][5] & ~x[0];
			partial_clause[4][6] 	= partial_clause_prev[4][6] & 1'b1;
			partial_clause[4][7] 	= partial_clause_prev[4][7] & ~x[15];
			partial_clause[4][8] 	= partial_clause_prev[4][8] & 1'b1;
			partial_clause[4][9] 	= partial_clause_prev[4][9] & 1'b1;
			partial_clause[4][10] 	= partial_clause_prev[4][10] & 1'b1;
			partial_clause[4][11] 	= partial_clause_prev[4][11] & 1'b1;
			partial_clause[4][12] 	= partial_clause_prev[4][12] & 1'b1;
			partial_clause[4][13] 	= partial_clause_prev[4][13] & 1'b1;
			partial_clause[4][14] 	= partial_clause_prev[4][14] & 1'b1;
			partial_clause[4][15] 	= partial_clause_prev[4][15] & 1'b1;
			partial_clause[4][16] 	= partial_clause_prev[4][16] & 1'b1;
			partial_clause[4][17] 	= partial_clause_prev[4][17] & 1'b1;
			partial_clause[4][18] 	= partial_clause_prev[4][18] & 1'b1;
			partial_clause[4][19] 	= partial_clause_prev[4][19] & 1'b1;
			partial_clause[4][20] 	= partial_clause_prev[4][20] & 1'b1;
			partial_clause[4][21] 	= partial_clause_prev[4][21] & 1'b1;
			partial_clause[4][22] 	= partial_clause_prev[4][22] & 1'b1;
			partial_clause[4][23] 	= partial_clause_prev[4][23] & 1'b1;
			partial_clause[4][24] 	= partial_clause_prev[4][24] & 1'b1;
			partial_clause[4][25] 	= partial_clause_prev[4][25] & ~x[12];
			partial_clause[4][26] 	= partial_clause_prev[4][26] & 1'b1;
			partial_clause[4][27] 	= partial_clause_prev[4][27] & 1'b1;
			partial_clause[4][28] 	= partial_clause_prev[4][28] & 1'b1;
			partial_clause[4][29] 	= partial_clause_prev[4][29] & 1'b1;
			partial_clause[4][30] 	= partial_clause_prev[4][30] & 1'b1;
			partial_clause[4][31] 	= partial_clause_prev[4][31] & 1'b1;
			partial_clause[4][32] 	= partial_clause_prev[4][32] & 1'b1;
			partial_clause[4][33] 	= partial_clause_prev[4][33] & ~x[1];
			partial_clause[4][34] 	= partial_clause_prev[4][34] & 1'b1;
			partial_clause[4][35] 	= partial_clause_prev[4][35] & 1'b1;
			partial_clause[4][36] 	= partial_clause_prev[4][36] & 1'b1;
			partial_clause[4][37] 	= partial_clause_prev[4][37] & 1'b1;
			partial_clause[4][38] 	= partial_clause_prev[4][38] & 1'b1;
			partial_clause[4][39] 	= partial_clause_prev[4][39] & 1'b1;
			partial_clause[4][40] 	= partial_clause_prev[4][40] & 1'b1;
			partial_clause[4][41] 	= partial_clause_prev[4][41] & 1'b1;
			partial_clause[4][42] 	= partial_clause_prev[4][42] & 1'b1;
			partial_clause[4][43] 	= partial_clause_prev[4][43] & 1'b1;
			partial_clause[4][44] 	= partial_clause_prev[4][44] & 1'b1;
			partial_clause[4][45] 	= partial_clause_prev[4][45] & 1'b1;
			partial_clause[4][46] 	= partial_clause_prev[4][46] & 1'b1;
			partial_clause[4][47] 	= partial_clause_prev[4][47] & 1'b1;
			partial_clause[4][48] 	= partial_clause_prev[4][48] & 1'b1;
			partial_clause[4][49] 	= partial_clause_prev[4][49] & ~x[5];
			partial_clause[4][50] 	= partial_clause_prev[4][50] & ~x[7];
			partial_clause[4][51] 	= partial_clause_prev[4][51] & ~x[13];
			partial_clause[4][52] 	= partial_clause_prev[4][52] & 1'b1;
			partial_clause[4][53] 	= partial_clause_prev[4][53] & 1'b1;
			partial_clause[4][54] 	= partial_clause_prev[4][54] & 1'b1;
			partial_clause[4][55] 	= partial_clause_prev[4][55] & 1'b1;
			partial_clause[4][56] 	= partial_clause_prev[4][56] & 1'b1;
			partial_clause[4][57] 	= partial_clause_prev[4][57] & 1'b1;
			partial_clause[4][58] 	= partial_clause_prev[4][58] & ~x[14];
			partial_clause[4][59] 	= partial_clause_prev[4][59] & 1'b1;
			partial_clause[4][60] 	= partial_clause_prev[4][60] & ~x[0];
			partial_clause[4][61] 	= partial_clause_prev[4][61] & ~x[1];
			partial_clause[4][62] 	= partial_clause_prev[4][62] & 1'b1;
			partial_clause[4][63] 	= partial_clause_prev[4][63] & ~x[11];
			partial_clause[4][64] 	= partial_clause_prev[4][64] & ~x[10];
			partial_clause[4][65] 	= partial_clause_prev[4][65] & 1'b1;
			partial_clause[4][66] 	= partial_clause_prev[4][66] & 1'b1;
			partial_clause[4][67] 	= partial_clause_prev[4][67] & 1'b1;
			partial_clause[4][68] 	= partial_clause_prev[4][68] & ~x[4];
			partial_clause[4][69] 	= partial_clause_prev[4][69] & 1'b1;
			partial_clause[4][70] 	= partial_clause_prev[4][70] & 1'b1;
			partial_clause[4][71] 	= partial_clause_prev[4][71] & 1'b1;
			partial_clause[4][72] 	= partial_clause_prev[4][72] & 1'b1;
			partial_clause[4][73] 	= partial_clause_prev[4][73] & ~x[0];
			partial_clause[4][74] 	= partial_clause_prev[4][74] & 1'b1;
			partial_clause[4][75] 	= partial_clause_prev[4][75] & 1'b1;
			partial_clause[4][76] 	= partial_clause_prev[4][76] & ~x[4];
			partial_clause[4][77] 	= partial_clause_prev[4][77] & 1'b1;
			partial_clause[4][78] 	= partial_clause_prev[4][78] & 1'b1;
			partial_clause[4][79] 	= partial_clause_prev[4][79] & ~x[13];
			partial_clause[4][80] 	= partial_clause_prev[4][80] & 1'b1;
			partial_clause[4][81] 	= partial_clause_prev[4][81] & 1'b1;
			partial_clause[4][82] 	= partial_clause_prev[4][82] & 1'b1;
			partial_clause[4][83] 	= partial_clause_prev[4][83] & 1'b1;
			partial_clause[4][84] 	= partial_clause_prev[4][84] & 1'b1;
			partial_clause[4][85] 	= partial_clause_prev[4][85] & 1'b1;
			partial_clause[4][86] 	= partial_clause_prev[4][86] & 1'b1;
			partial_clause[4][87] 	= partial_clause_prev[4][87] & 1'b1;
			partial_clause[4][88] 	= partial_clause_prev[4][88] & 1'b1;
			partial_clause[4][89] 	= partial_clause_prev[4][89] & 1'b1;
			partial_clause[4][90] 	= partial_clause_prev[4][90] & 1'b1;
			partial_clause[4][91] 	= partial_clause_prev[4][91] & 1'b1;
			partial_clause[4][92] 	= partial_clause_prev[4][92] & 1'b1;
			partial_clause[4][93] 	= partial_clause_prev[4][93] & 1'b1;
			partial_clause[4][94] 	= partial_clause_prev[4][94] & 1'b1;
			partial_clause[4][95] 	= partial_clause_prev[4][95] & 1'b1;
			partial_clause[4][96] 	= partial_clause_prev[4][96] & 1'b1;
			partial_clause[4][97] 	= partial_clause_prev[4][97] & ~x[14];
			partial_clause[4][98] 	= partial_clause_prev[4][98] & 1'b1;
			partial_clause[4][99] 	= partial_clause_prev[4][99] & 1'b1;
			// Class 5
			partial_clause[5][0] 	= partial_clause_prev[5][0] & 1'b1;
			partial_clause[5][1] 	= partial_clause_prev[5][1] & 1'b1;
			partial_clause[5][2] 	= partial_clause_prev[5][2] & 1'b1;
			partial_clause[5][3] 	= partial_clause_prev[5][3] & 1'b1;
			partial_clause[5][4] 	= partial_clause_prev[5][4] & 1'b1;
			partial_clause[5][5] 	= partial_clause_prev[5][5] & 1'b1;
			partial_clause[5][6] 	= partial_clause_prev[5][6] & 1'b1;
			partial_clause[5][7] 	= partial_clause_prev[5][7] & 1'b1;
			partial_clause[5][8] 	= partial_clause_prev[5][8] & ~x[0];
			partial_clause[5][9] 	= partial_clause_prev[5][9] & 1'b1;
			partial_clause[5][10] 	= partial_clause_prev[5][10] & 1'b1;
			partial_clause[5][11] 	= partial_clause_prev[5][11] & 1'b1;
			partial_clause[5][12] 	= partial_clause_prev[5][12] & 1'b1;
			partial_clause[5][13] 	= partial_clause_prev[5][13] & 1'b1;
			partial_clause[5][14] 	= partial_clause_prev[5][14] & 1'b1;
			partial_clause[5][15] 	= partial_clause_prev[5][15] & 1'b1;
			partial_clause[5][16] 	= partial_clause_prev[5][16] & 1'b1;
			partial_clause[5][17] 	= partial_clause_prev[5][17] & 1'b1;
			partial_clause[5][18] 	= partial_clause_prev[5][18] & 1'b1;
			partial_clause[5][19] 	= partial_clause_prev[5][19] & 1'b1;
			partial_clause[5][20] 	= partial_clause_prev[5][20] & 1'b1;
			partial_clause[5][21] 	= partial_clause_prev[5][21] & 1'b1;
			partial_clause[5][22] 	= partial_clause_prev[5][22] & 1'b1;
			partial_clause[5][23] 	= partial_clause_prev[5][23] & 1'b1;
			partial_clause[5][24] 	= partial_clause_prev[5][24] & 1'b1;
			partial_clause[5][25] 	= partial_clause_prev[5][25] & 1'b1;
			partial_clause[5][26] 	= partial_clause_prev[5][26] & 1'b1;
			partial_clause[5][27] 	= partial_clause_prev[5][27] & 1'b1;
			partial_clause[5][28] 	= partial_clause_prev[5][28] & 1'b1;
			partial_clause[5][29] 	= partial_clause_prev[5][29] & 1'b1;
			partial_clause[5][30] 	= partial_clause_prev[5][30] & 1'b1;
			partial_clause[5][31] 	= partial_clause_prev[5][31] & 1'b1;
			partial_clause[5][32] 	= partial_clause_prev[5][32] & 1'b1;
			partial_clause[5][33] 	= partial_clause_prev[5][33] & 1'b1;
			partial_clause[5][34] 	= partial_clause_prev[5][34] & 1'b1;
			partial_clause[5][35] 	= partial_clause_prev[5][35] & 1'b1;
			partial_clause[5][36] 	= partial_clause_prev[5][36] & 1'b1;
			partial_clause[5][37] 	= partial_clause_prev[5][37] & 1'b1;
			partial_clause[5][38] 	= partial_clause_prev[5][38] & 1'b1;
			partial_clause[5][39] 	= partial_clause_prev[5][39] & 1'b1;
			partial_clause[5][40] 	= partial_clause_prev[5][40] & 1'b1;
			partial_clause[5][41] 	= partial_clause_prev[5][41] & 1'b1;
			partial_clause[5][42] 	= partial_clause_prev[5][42] & ~x[12];
			partial_clause[5][43] 	= partial_clause_prev[5][43] & 1'b1;
			partial_clause[5][44] 	= partial_clause_prev[5][44] & 1'b1;
			partial_clause[5][45] 	= partial_clause_prev[5][45] & 1'b1;
			partial_clause[5][46] 	= partial_clause_prev[5][46] & 1'b1;
			partial_clause[5][47] 	= partial_clause_prev[5][47] & 1'b1;
			partial_clause[5][48] 	= partial_clause_prev[5][48] & 1'b1;
			partial_clause[5][49] 	= partial_clause_prev[5][49] & 1'b1;
			partial_clause[5][50] 	= partial_clause_prev[5][50] & 1'b1;
			partial_clause[5][51] 	= partial_clause_prev[5][51] & 1'b1;
			partial_clause[5][52] 	= partial_clause_prev[5][52] & 1'b1;
			partial_clause[5][53] 	= partial_clause_prev[5][53] & 1'b1;
			partial_clause[5][54] 	= partial_clause_prev[5][54] & 1'b1;
			partial_clause[5][55] 	= partial_clause_prev[5][55] & 1'b1;
			partial_clause[5][56] 	= partial_clause_prev[5][56] & 1'b1;
			partial_clause[5][57] 	= partial_clause_prev[5][57] & 1'b1;
			partial_clause[5][58] 	= partial_clause_prev[5][58] & 1'b1;
			partial_clause[5][59] 	= partial_clause_prev[5][59] & 1'b1;
			partial_clause[5][60] 	= partial_clause_prev[5][60] & 1'b1;
			partial_clause[5][61] 	= partial_clause_prev[5][61] & 1'b1;
			partial_clause[5][62] 	= partial_clause_prev[5][62] & 1'b1;
			partial_clause[5][63] 	= partial_clause_prev[5][63] & 1'b1;
			partial_clause[5][64] 	= partial_clause_prev[5][64] & ~x[11];
			partial_clause[5][65] 	= partial_clause_prev[5][65] & 1'b1;
			partial_clause[5][66] 	= partial_clause_prev[5][66] & ~x[11];
			partial_clause[5][67] 	= partial_clause_prev[5][67] & 1'b1;
			partial_clause[5][68] 	= partial_clause_prev[5][68] & 1'b1;
			partial_clause[5][69] 	= partial_clause_prev[5][69] & 1'b1;
			partial_clause[5][70] 	= partial_clause_prev[5][70] & 1'b1;
			partial_clause[5][71] 	= partial_clause_prev[5][71] & 1'b1;
			partial_clause[5][72] 	= partial_clause_prev[5][72] & 1'b1;
			partial_clause[5][73] 	= partial_clause_prev[5][73] & 1'b1;
			partial_clause[5][74] 	= partial_clause_prev[5][74] & ~x[6];
			partial_clause[5][75] 	= partial_clause_prev[5][75] & 1'b1;
			partial_clause[5][76] 	= partial_clause_prev[5][76] & 1'b1;
			partial_clause[5][77] 	= partial_clause_prev[5][77] & ~x[6];
			partial_clause[5][78] 	= partial_clause_prev[5][78] & ~x[10];
			partial_clause[5][79] 	= partial_clause_prev[5][79] & 1'b1;
			partial_clause[5][80] 	= partial_clause_prev[5][80] & 1'b1;
			partial_clause[5][81] 	= partial_clause_prev[5][81] & 1'b1;
			partial_clause[5][82] 	= partial_clause_prev[5][82] & 1'b1;
			partial_clause[5][83] 	= partial_clause_prev[5][83] & 1'b1;
			partial_clause[5][84] 	= partial_clause_prev[5][84] & 1'b1;
			partial_clause[5][85] 	= partial_clause_prev[5][85] & 1'b1;
			partial_clause[5][86] 	= partial_clause_prev[5][86] & 1'b1;
			partial_clause[5][87] 	= partial_clause_prev[5][87] & 1'b1;
			partial_clause[5][88] 	= partial_clause_prev[5][88] & 1'b1;
			partial_clause[5][89] 	= partial_clause_prev[5][89] & 1'b1;
			partial_clause[5][90] 	= partial_clause_prev[5][90] & ~x[13];
			partial_clause[5][91] 	= partial_clause_prev[5][91] & 1'b1;
			partial_clause[5][92] 	= partial_clause_prev[5][92] & 1'b1;
			partial_clause[5][93] 	= partial_clause_prev[5][93] & 1'b1;
			partial_clause[5][94] 	= partial_clause_prev[5][94] & 1'b1;
			partial_clause[5][95] 	= partial_clause_prev[5][95] & 1'b1;
			partial_clause[5][96] 	= partial_clause_prev[5][96] & 1'b1;
			partial_clause[5][97] 	= partial_clause_prev[5][97] & 1'b1;
			partial_clause[5][98] 	= partial_clause_prev[5][98] & 1'b1;
			partial_clause[5][99] 	= partial_clause_prev[5][99] & 1'b1;
			// Class 6
			partial_clause[6][0] 	= partial_clause_prev[6][0] & 1'b1;
			partial_clause[6][1] 	= partial_clause_prev[6][1] & ~x[0];
			partial_clause[6][2] 	= partial_clause_prev[6][2] & 1'b1;
			partial_clause[6][3] 	= partial_clause_prev[6][3] & 1'b1;
			partial_clause[6][4] 	= partial_clause_prev[6][4] & ~x[7];
			partial_clause[6][5] 	= partial_clause_prev[6][5] & 1'b1;
			partial_clause[6][6] 	= partial_clause_prev[6][6] & 1'b1;
			partial_clause[6][7] 	= partial_clause_prev[6][7] & 1'b1;
			partial_clause[6][8] 	= partial_clause_prev[6][8] & 1'b1;
			partial_clause[6][9] 	= partial_clause_prev[6][9] & 1'b1;
			partial_clause[6][10] 	= partial_clause_prev[6][10] & 1'b1;
			partial_clause[6][11] 	= partial_clause_prev[6][11] & 1'b1;
			partial_clause[6][12] 	= partial_clause_prev[6][12] & 1'b1;
			partial_clause[6][13] 	= partial_clause_prev[6][13] & 1'b1;
			partial_clause[6][14] 	= partial_clause_prev[6][14] & 1'b1;
			partial_clause[6][15] 	= partial_clause_prev[6][15] & 1'b1;
			partial_clause[6][16] 	= partial_clause_prev[6][16] & 1'b1;
			partial_clause[6][17] 	= partial_clause_prev[6][17] & 1'b1;
			partial_clause[6][18] 	= partial_clause_prev[6][18] & 1'b1;
			partial_clause[6][19] 	= partial_clause_prev[6][19] & 1'b1;
			partial_clause[6][20] 	= partial_clause_prev[6][20] & 1'b1;
			partial_clause[6][21] 	= partial_clause_prev[6][21] & 1'b1;
			partial_clause[6][22] 	= partial_clause_prev[6][22] & 1'b1;
			partial_clause[6][23] 	= partial_clause_prev[6][23] & 1'b1;
			partial_clause[6][24] 	= partial_clause_prev[6][24] & 1'b1;
			partial_clause[6][25] 	= partial_clause_prev[6][25] & 1'b1;
			partial_clause[6][26] 	= partial_clause_prev[6][26] & 1'b1;
			partial_clause[6][27] 	= partial_clause_prev[6][27] & 1'b1;
			partial_clause[6][28] 	= partial_clause_prev[6][28] & 1'b1;
			partial_clause[6][29] 	= partial_clause_prev[6][29] & 1'b1;
			partial_clause[6][30] 	= partial_clause_prev[6][30] & 1'b1;
			partial_clause[6][31] 	= partial_clause_prev[6][31] & 1'b1;
			partial_clause[6][32] 	= partial_clause_prev[6][32] & 1'b1;
			partial_clause[6][33] 	= partial_clause_prev[6][33] & 1'b1;
			partial_clause[6][34] 	= partial_clause_prev[6][34] & 1'b1;
			partial_clause[6][35] 	= partial_clause_prev[6][35] & 1'b1;
			partial_clause[6][36] 	= partial_clause_prev[6][36] & 1'b1;
			partial_clause[6][37] 	= partial_clause_prev[6][37] & 1'b1;
			partial_clause[6][38] 	= partial_clause_prev[6][38] & 1'b1;
			partial_clause[6][39] 	= partial_clause_prev[6][39] & 1'b1;
			partial_clause[6][40] 	= partial_clause_prev[6][40] & 1'b1;
			partial_clause[6][41] 	= partial_clause_prev[6][41] & 1'b1;
			partial_clause[6][42] 	= partial_clause_prev[6][42] & 1'b1;
			partial_clause[6][43] 	= partial_clause_prev[6][43] & 1'b1;
			partial_clause[6][44] 	= partial_clause_prev[6][44] & 1'b1;
			partial_clause[6][45] 	= partial_clause_prev[6][45] & 1'b1;
			partial_clause[6][46] 	= partial_clause_prev[6][46] & 1'b1;
			partial_clause[6][47] 	= partial_clause_prev[6][47] & 1'b1;
			partial_clause[6][48] 	= partial_clause_prev[6][48] & 1'b1;
			partial_clause[6][49] 	= partial_clause_prev[6][49] & 1'b1;
			partial_clause[6][50] 	= partial_clause_prev[6][50] & 1'b1;
			partial_clause[6][51] 	= partial_clause_prev[6][51] & 1'b1;
			partial_clause[6][52] 	= partial_clause_prev[6][52] & 1'b1;
			partial_clause[6][53] 	= partial_clause_prev[6][53] & 1'b1;
			partial_clause[6][54] 	= partial_clause_prev[6][54] & 1'b1;
			partial_clause[6][55] 	= partial_clause_prev[6][55] & 1'b1;
			partial_clause[6][56] 	= partial_clause_prev[6][56] & 1'b1;
			partial_clause[6][57] 	= partial_clause_prev[6][57] & 1'b1;
			partial_clause[6][58] 	= partial_clause_prev[6][58] & 1'b1;
			partial_clause[6][59] 	= partial_clause_prev[6][59] & 1'b1;
			partial_clause[6][60] 	= partial_clause_prev[6][60] & 1'b1;
			partial_clause[6][61] 	= partial_clause_prev[6][61] & 1'b1;
			partial_clause[6][62] 	= partial_clause_prev[6][62] & 1'b1;
			partial_clause[6][63] 	= partial_clause_prev[6][63] & 1'b1;
			partial_clause[6][64] 	= partial_clause_prev[6][64] & 1'b1;
			partial_clause[6][65] 	= partial_clause_prev[6][65] & 1'b1;
			partial_clause[6][66] 	= partial_clause_prev[6][66] & 1'b1;
			partial_clause[6][67] 	= partial_clause_prev[6][67] & 1'b1;
			partial_clause[6][68] 	= partial_clause_prev[6][68] & 1'b1;
			partial_clause[6][69] 	= partial_clause_prev[6][69] & 1'b1;
			partial_clause[6][70] 	= partial_clause_prev[6][70] & 1'b1;
			partial_clause[6][71] 	= partial_clause_prev[6][71] & 1'b1;
			partial_clause[6][72] 	= partial_clause_prev[6][72] & 1'b1;
			partial_clause[6][73] 	= partial_clause_prev[6][73] & 1'b1;
			partial_clause[6][74] 	= partial_clause_prev[6][74] & ~x[2];
			partial_clause[6][75] 	= partial_clause_prev[6][75] & 1'b1;
			partial_clause[6][76] 	= partial_clause_prev[6][76] & 1'b1;
			partial_clause[6][77] 	= partial_clause_prev[6][77] & 1'b1;
			partial_clause[6][78] 	= partial_clause_prev[6][78] & 1'b1;
			partial_clause[6][79] 	= partial_clause_prev[6][79] & 1'b1;
			partial_clause[6][80] 	= partial_clause_prev[6][80] & 1'b1;
			partial_clause[6][81] 	= partial_clause_prev[6][81] & 1'b1;
			partial_clause[6][82] 	= partial_clause_prev[6][82] & 1'b1;
			partial_clause[6][83] 	= partial_clause_prev[6][83] & 1'b1;
			partial_clause[6][84] 	= partial_clause_prev[6][84] & 1'b1;
			partial_clause[6][85] 	= partial_clause_prev[6][85] & 1'b1;
			partial_clause[6][86] 	= partial_clause_prev[6][86] & 1'b1;
			partial_clause[6][87] 	= partial_clause_prev[6][87] & ~x[6];
			partial_clause[6][88] 	= partial_clause_prev[6][88] & 1'b1;
			partial_clause[6][89] 	= partial_clause_prev[6][89] & 1'b1;
			partial_clause[6][90] 	= partial_clause_prev[6][90] & 1'b1;
			partial_clause[6][91] 	= partial_clause_prev[6][91] & ~x[5];
			partial_clause[6][92] 	= partial_clause_prev[6][92] & 1'b1;
			partial_clause[6][93] 	= partial_clause_prev[6][93] & 1'b1;
			partial_clause[6][94] 	= partial_clause_prev[6][94] & 1'b1;
			partial_clause[6][95] 	= partial_clause_prev[6][95] & ~x[10];
			partial_clause[6][96] 	= partial_clause_prev[6][96] & ~x[4];
			partial_clause[6][97] 	= partial_clause_prev[6][97] & 1'b1;
			partial_clause[6][98] 	= partial_clause_prev[6][98] & 1'b1;
			partial_clause[6][99] 	= partial_clause_prev[6][99] & 1'b1;
			// Class 7
			partial_clause[7][0] 	= partial_clause_prev[7][0] & 1'b1;
			partial_clause[7][1] 	= partial_clause_prev[7][1] & 1'b1;
			partial_clause[7][2] 	= partial_clause_prev[7][2] & 1'b1;
			partial_clause[7][3] 	= partial_clause_prev[7][3] & 1'b1;
			partial_clause[7][4] 	= partial_clause_prev[7][4] & 1'b1;
			partial_clause[7][5] 	= partial_clause_prev[7][5] & 1'b1;
			partial_clause[7][6] 	= partial_clause_prev[7][6] & 1'b1;
			partial_clause[7][7] 	= partial_clause_prev[7][7] & 1'b1;
			partial_clause[7][8] 	= partial_clause_prev[7][8] & 1'b1;
			partial_clause[7][9] 	= partial_clause_prev[7][9] & 1'b1;
			partial_clause[7][10] 	= partial_clause_prev[7][10] & 1'b1;
			partial_clause[7][11] 	= partial_clause_prev[7][11] & 1'b1;
			partial_clause[7][12] 	= partial_clause_prev[7][12] & 1'b1;
			partial_clause[7][13] 	= partial_clause_prev[7][13] & 1'b1;
			partial_clause[7][14] 	= partial_clause_prev[7][14] & 1'b1;
			partial_clause[7][15] 	= partial_clause_prev[7][15] & 1'b1;
			partial_clause[7][16] 	= partial_clause_prev[7][16] & 1'b1;
			partial_clause[7][17] 	= partial_clause_prev[7][17] & 1'b1;
			partial_clause[7][18] 	= partial_clause_prev[7][18] & 1'b1;
			partial_clause[7][19] 	= partial_clause_prev[7][19] & 1'b1;
			partial_clause[7][20] 	= partial_clause_prev[7][20] & 1'b1;
			partial_clause[7][21] 	= partial_clause_prev[7][21] & 1'b1;
			partial_clause[7][22] 	= partial_clause_prev[7][22] & 1'b1;
			partial_clause[7][23] 	= partial_clause_prev[7][23] & 1'b1;
			partial_clause[7][24] 	= partial_clause_prev[7][24] & 1'b1;
			partial_clause[7][25] 	= partial_clause_prev[7][25] & 1'b1;
			partial_clause[7][26] 	= partial_clause_prev[7][26] & 1'b1;
			partial_clause[7][27] 	= partial_clause_prev[7][27] & 1'b1;
			partial_clause[7][28] 	= partial_clause_prev[7][28] & 1'b1;
			partial_clause[7][29] 	= partial_clause_prev[7][29] & 1'b1;
			partial_clause[7][30] 	= partial_clause_prev[7][30] & 1'b1;
			partial_clause[7][31] 	= partial_clause_prev[7][31] & 1'b1;
			partial_clause[7][32] 	= partial_clause_prev[7][32] & 1'b1;
			partial_clause[7][33] 	= partial_clause_prev[7][33] & 1'b1;
			partial_clause[7][34] 	= partial_clause_prev[7][34] & 1'b1;
			partial_clause[7][35] 	= partial_clause_prev[7][35] & 1'b1;
			partial_clause[7][36] 	= partial_clause_prev[7][36] & 1'b1;
			partial_clause[7][37] 	= partial_clause_prev[7][37] & 1'b1;
			partial_clause[7][38] 	= partial_clause_prev[7][38] & ~x[14];
			partial_clause[7][39] 	= partial_clause_prev[7][39] & 1'b1;
			partial_clause[7][40] 	= partial_clause_prev[7][40] & 1'b1;
			partial_clause[7][41] 	= partial_clause_prev[7][41] & 1'b1;
			partial_clause[7][42] 	= partial_clause_prev[7][42] & 1'b1;
			partial_clause[7][43] 	= partial_clause_prev[7][43] & 1'b1;
			partial_clause[7][44] 	= partial_clause_prev[7][44] & 1'b1;
			partial_clause[7][45] 	= partial_clause_prev[7][45] & 1'b1;
			partial_clause[7][46] 	= partial_clause_prev[7][46] & 1'b1;
			partial_clause[7][47] 	= partial_clause_prev[7][47] & 1'b1;
			partial_clause[7][48] 	= partial_clause_prev[7][48] & 1'b1;
			partial_clause[7][49] 	= partial_clause_prev[7][49] & 1'b1;
			partial_clause[7][50] 	= partial_clause_prev[7][50] & 1'b1;
			partial_clause[7][51] 	= partial_clause_prev[7][51] & 1'b1;
			partial_clause[7][52] 	= partial_clause_prev[7][52] & ~x[2];
			partial_clause[7][53] 	= partial_clause_prev[7][53] & 1'b1;
			partial_clause[7][54] 	= partial_clause_prev[7][54] & ~x[8];
			partial_clause[7][55] 	= partial_clause_prev[7][55] & 1'b1;
			partial_clause[7][56] 	= partial_clause_prev[7][56] & 1'b1;
			partial_clause[7][57] 	= partial_clause_prev[7][57] & 1'b1;
			partial_clause[7][58] 	= partial_clause_prev[7][58] & ~x[0];
			partial_clause[7][59] 	= partial_clause_prev[7][59] & 1'b1;
			partial_clause[7][60] 	= partial_clause_prev[7][60] & 1'b1;
			partial_clause[7][61] 	= partial_clause_prev[7][61] & 1'b1;
			partial_clause[7][62] 	= partial_clause_prev[7][62] & 1'b1;
			partial_clause[7][63] 	= partial_clause_prev[7][63] & 1'b1;
			partial_clause[7][64] 	= partial_clause_prev[7][64] & 1'b1;
			partial_clause[7][65] 	= partial_clause_prev[7][65] & 1'b1;
			partial_clause[7][66] 	= partial_clause_prev[7][66] & ~x[15];
			partial_clause[7][67] 	= partial_clause_prev[7][67] & 1'b1;
			partial_clause[7][68] 	= partial_clause_prev[7][68] & 1'b1;
			partial_clause[7][69] 	= partial_clause_prev[7][69] & 1'b1;
			partial_clause[7][70] 	= partial_clause_prev[7][70] & 1'b1;
			partial_clause[7][71] 	= partial_clause_prev[7][71] & 1'b1;
			partial_clause[7][72] 	= partial_clause_prev[7][72] & 1'b1;
			partial_clause[7][73] 	= partial_clause_prev[7][73] & 1'b1;
			partial_clause[7][74] 	= partial_clause_prev[7][74] & 1'b1;
			partial_clause[7][75] 	= partial_clause_prev[7][75] & ~x[7];
			partial_clause[7][76] 	= partial_clause_prev[7][76] & 1'b1;
			partial_clause[7][77] 	= partial_clause_prev[7][77] & 1'b1;
			partial_clause[7][78] 	= partial_clause_prev[7][78] & ~x[2];
			partial_clause[7][79] 	= partial_clause_prev[7][79] & 1'b1;
			partial_clause[7][80] 	= partial_clause_prev[7][80] & 1'b1;
			partial_clause[7][81] 	= partial_clause_prev[7][81] & 1'b1;
			partial_clause[7][82] 	= partial_clause_prev[7][82] & ~x[6];
			partial_clause[7][83] 	= partial_clause_prev[7][83] & 1'b1;
			partial_clause[7][84] 	= partial_clause_prev[7][84] & 1'b1;
			partial_clause[7][85] 	= partial_clause_prev[7][85] & 1'b1;
			partial_clause[7][86] 	= partial_clause_prev[7][86] & 1'b1;
			partial_clause[7][87] 	= partial_clause_prev[7][87] & 1'b1;
			partial_clause[7][88] 	= partial_clause_prev[7][88] & ~x[2];
			partial_clause[7][89] 	= partial_clause_prev[7][89] & 1'b1;
			partial_clause[7][90] 	= partial_clause_prev[7][90] & 1'b1;
			partial_clause[7][91] 	= partial_clause_prev[7][91] & 1'b1;
			partial_clause[7][92] 	= partial_clause_prev[7][92] & 1'b1;
			partial_clause[7][93] 	= partial_clause_prev[7][93] & 1'b1;
			partial_clause[7][94] 	= partial_clause_prev[7][94] & 1'b1;
			partial_clause[7][95] 	= partial_clause_prev[7][95] & ~x[5];
			partial_clause[7][96] 	= partial_clause_prev[7][96] & 1'b1;
			partial_clause[7][97] 	= partial_clause_prev[7][97] & 1'b1;
			partial_clause[7][98] 	= partial_clause_prev[7][98] & 1'b1;
			partial_clause[7][99] 	= partial_clause_prev[7][99] & 1'b1;
			// Class 8
			partial_clause[8][0] 	= partial_clause_prev[8][0] & ~x[9];
			partial_clause[8][1] 	= partial_clause_prev[8][1] & ~x[0];
			partial_clause[8][2] 	= partial_clause_prev[8][2] & 1'b1;
			partial_clause[8][3] 	= partial_clause_prev[8][3] & 1'b1;
			partial_clause[8][4] 	= partial_clause_prev[8][4] & 1'b1;
			partial_clause[8][5] 	= partial_clause_prev[8][5] & 1'b1;
			partial_clause[8][6] 	= partial_clause_prev[8][6] & 1'b1;
			partial_clause[8][7] 	= partial_clause_prev[8][7] & 1'b1;
			partial_clause[8][8] 	= partial_clause_prev[8][8] & 1'b1;
			partial_clause[8][9] 	= partial_clause_prev[8][9] & 1'b1;
			partial_clause[8][10] 	= partial_clause_prev[8][10] & 1'b1;
			partial_clause[8][11] 	= partial_clause_prev[8][11] & 1'b1;
			partial_clause[8][12] 	= partial_clause_prev[8][12] & 1'b1;
			partial_clause[8][13] 	= partial_clause_prev[8][13] & 1'b1;
			partial_clause[8][14] 	= partial_clause_prev[8][14] & 1'b1;
			partial_clause[8][15] 	= partial_clause_prev[8][15] & 1'b1;
			partial_clause[8][16] 	= partial_clause_prev[8][16] & 1'b1;
			partial_clause[8][17] 	= partial_clause_prev[8][17] & 1'b1;
			partial_clause[8][18] 	= partial_clause_prev[8][18] & 1'b1;
			partial_clause[8][19] 	= partial_clause_prev[8][19] & 1'b1;
			partial_clause[8][20] 	= partial_clause_prev[8][20] & 1'b1;
			partial_clause[8][21] 	= partial_clause_prev[8][21] & ~x[1];
			partial_clause[8][22] 	= partial_clause_prev[8][22] & 1'b1;
			partial_clause[8][23] 	= partial_clause_prev[8][23] & 1'b1;
			partial_clause[8][24] 	= partial_clause_prev[8][24] & ~x[14];
			partial_clause[8][25] 	= partial_clause_prev[8][25] & 1'b1;
			partial_clause[8][26] 	= partial_clause_prev[8][26] & 1'b1;
			partial_clause[8][27] 	= partial_clause_prev[8][27] & 1'b1;
			partial_clause[8][28] 	= partial_clause_prev[8][28] & 1'b1;
			partial_clause[8][29] 	= partial_clause_prev[8][29] & 1'b1;
			partial_clause[8][30] 	= partial_clause_prev[8][30] & 1'b1;
			partial_clause[8][31] 	= partial_clause_prev[8][31] & 1'b1;
			partial_clause[8][32] 	= partial_clause_prev[8][32] & ~x[1];
			partial_clause[8][33] 	= partial_clause_prev[8][33] & 1'b1;
			partial_clause[8][34] 	= partial_clause_prev[8][34] & 1'b1;
			partial_clause[8][35] 	= partial_clause_prev[8][35] & 1'b1;
			partial_clause[8][36] 	= partial_clause_prev[8][36] & 1'b1;
			partial_clause[8][37] 	= partial_clause_prev[8][37] & 1'b1;
			partial_clause[8][38] 	= partial_clause_prev[8][38] & 1'b1;
			partial_clause[8][39] 	= partial_clause_prev[8][39] & 1'b1;
			partial_clause[8][40] 	= partial_clause_prev[8][40] & 1'b1;
			partial_clause[8][41] 	= partial_clause_prev[8][41] & 1'b1;
			partial_clause[8][42] 	= partial_clause_prev[8][42] & 1'b1;
			partial_clause[8][43] 	= partial_clause_prev[8][43] & 1'b1;
			partial_clause[8][44] 	= partial_clause_prev[8][44] & ~x[3];
			partial_clause[8][45] 	= partial_clause_prev[8][45] & 1'b1;
			partial_clause[8][46] 	= partial_clause_prev[8][46] & ~x[7] & ~x[9];
			partial_clause[8][47] 	= partial_clause_prev[8][47] & 1'b1;
			partial_clause[8][48] 	= partial_clause_prev[8][48] & 1'b1;
			partial_clause[8][49] 	= partial_clause_prev[8][49] & 1'b1;
			partial_clause[8][50] 	= partial_clause_prev[8][50] & ~x[7];
			partial_clause[8][51] 	= partial_clause_prev[8][51] & ~x[11];
			partial_clause[8][52] 	= partial_clause_prev[8][52] & 1'b1;
			partial_clause[8][53] 	= partial_clause_prev[8][53] & ~x[7];
			partial_clause[8][54] 	= partial_clause_prev[8][54] & ~x[10];
			partial_clause[8][55] 	= partial_clause_prev[8][55] & 1'b1;
			partial_clause[8][56] 	= partial_clause_prev[8][56] & 1'b1;
			partial_clause[8][57] 	= partial_clause_prev[8][57] & 1'b1;
			partial_clause[8][58] 	= partial_clause_prev[8][58] & 1'b1;
			partial_clause[8][59] 	= partial_clause_prev[8][59] & 1'b1;
			partial_clause[8][60] 	= partial_clause_prev[8][60] & 1'b1;
			partial_clause[8][61] 	= partial_clause_prev[8][61] & 1'b1;
			partial_clause[8][62] 	= partial_clause_prev[8][62] & ~x[14];
			partial_clause[8][63] 	= partial_clause_prev[8][63] & 1'b1;
			partial_clause[8][64] 	= partial_clause_prev[8][64] & 1'b1;
			partial_clause[8][65] 	= partial_clause_prev[8][65] & 1'b1;
			partial_clause[8][66] 	= partial_clause_prev[8][66] & 1'b1;
			partial_clause[8][67] 	= partial_clause_prev[8][67] & 1'b1;
			partial_clause[8][68] 	= partial_clause_prev[8][68] & 1'b1;
			partial_clause[8][69] 	= partial_clause_prev[8][69] & 1'b1;
			partial_clause[8][70] 	= partial_clause_prev[8][70] & 1'b1;
			partial_clause[8][71] 	= partial_clause_prev[8][71] & 1'b1;
			partial_clause[8][72] 	= partial_clause_prev[8][72] & 1'b1;
			partial_clause[8][73] 	= partial_clause_prev[8][73] & 1'b1;
			partial_clause[8][74] 	= partial_clause_prev[8][74] & 1'b1;
			partial_clause[8][75] 	= partial_clause_prev[8][75] & 1'b1;
			partial_clause[8][76] 	= partial_clause_prev[8][76] & 1'b1;
			partial_clause[8][77] 	= partial_clause_prev[8][77] & 1'b1;
			partial_clause[8][78] 	= partial_clause_prev[8][78] & 1'b1;
			partial_clause[8][79] 	= partial_clause_prev[8][79] & 1'b1;
			partial_clause[8][80] 	= partial_clause_prev[8][80] & 1'b1;
			partial_clause[8][81] 	= partial_clause_prev[8][81] & 1'b1;
			partial_clause[8][82] 	= partial_clause_prev[8][82] & 1'b1;
			partial_clause[8][83] 	= partial_clause_prev[8][83] & 1'b1;
			partial_clause[8][84] 	= partial_clause_prev[8][84] & ~x[3];
			partial_clause[8][85] 	= partial_clause_prev[8][85] & ~x[13];
			partial_clause[8][86] 	= partial_clause_prev[8][86] & ~x[3] & ~x[15];
			partial_clause[8][87] 	= partial_clause_prev[8][87] & 1'b1;
			partial_clause[8][88] 	= partial_clause_prev[8][88] & 1'b1;
			partial_clause[8][89] 	= partial_clause_prev[8][89] & ~x[8];
			partial_clause[8][90] 	= partial_clause_prev[8][90] & ~x[6];
			partial_clause[8][91] 	= partial_clause_prev[8][91] & 1'b1;
			partial_clause[8][92] 	= partial_clause_prev[8][92] & 1'b1;
			partial_clause[8][93] 	= partial_clause_prev[8][93] & 1'b1;
			partial_clause[8][94] 	= partial_clause_prev[8][94] & ~x[4];
			partial_clause[8][95] 	= partial_clause_prev[8][95] & ~x[5];
			partial_clause[8][96] 	= partial_clause_prev[8][96] & ~x[8];
			partial_clause[8][97] 	= partial_clause_prev[8][97] & 1'b1;
			partial_clause[8][98] 	= partial_clause_prev[8][98] & 1'b1;
			partial_clause[8][99] 	= partial_clause_prev[8][99] & 1'b1;
			// Class 9
			partial_clause[9][0] 	= partial_clause_prev[9][0] & 1'b1;
			partial_clause[9][1] 	= partial_clause_prev[9][1] & 1'b1;
			partial_clause[9][2] 	= partial_clause_prev[9][2] & 1'b1;
			partial_clause[9][3] 	= partial_clause_prev[9][3] & 1'b1;
			partial_clause[9][4] 	= partial_clause_prev[9][4] & 1'b1;
			partial_clause[9][5] 	= partial_clause_prev[9][5] & 1'b1;
			partial_clause[9][6] 	= partial_clause_prev[9][6] & 1'b1;
			partial_clause[9][7] 	= partial_clause_prev[9][7] & 1'b1;
			partial_clause[9][8] 	= partial_clause_prev[9][8] & 1'b1;
			partial_clause[9][9] 	= partial_clause_prev[9][9] & 1'b1;
			partial_clause[9][10] 	= partial_clause_prev[9][10] & 1'b1;
			partial_clause[9][11] 	= partial_clause_prev[9][11] & 1'b1;
			partial_clause[9][12] 	= partial_clause_prev[9][12] & 1'b1;
			partial_clause[9][13] 	= partial_clause_prev[9][13] & 1'b1;
			partial_clause[9][14] 	= partial_clause_prev[9][14] & 1'b1;
			partial_clause[9][15] 	= partial_clause_prev[9][15] & 1'b1;
			partial_clause[9][16] 	= partial_clause_prev[9][16] & 1'b1;
			partial_clause[9][17] 	= partial_clause_prev[9][17] & ~x[8];
			partial_clause[9][18] 	= partial_clause_prev[9][18] & 1'b1;
			partial_clause[9][19] 	= partial_clause_prev[9][19] & 1'b1;
			partial_clause[9][20] 	= partial_clause_prev[9][20] & 1'b1;
			partial_clause[9][21] 	= partial_clause_prev[9][21] & ~x[0];
			partial_clause[9][22] 	= partial_clause_prev[9][22] & 1'b1;
			partial_clause[9][23] 	= partial_clause_prev[9][23] & 1'b1;
			partial_clause[9][24] 	= partial_clause_prev[9][24] & 1'b1;
			partial_clause[9][25] 	= partial_clause_prev[9][25] & 1'b1;
			partial_clause[9][26] 	= partial_clause_prev[9][26] & 1'b1;
			partial_clause[9][27] 	= partial_clause_prev[9][27] & 1'b1;
			partial_clause[9][28] 	= partial_clause_prev[9][28] & 1'b1;
			partial_clause[9][29] 	= partial_clause_prev[9][29] & 1'b1;
			partial_clause[9][30] 	= partial_clause_prev[9][30] & 1'b1;
			partial_clause[9][31] 	= partial_clause_prev[9][31] & 1'b1;
			partial_clause[9][32] 	= partial_clause_prev[9][32] & 1'b1;
			partial_clause[9][33] 	= partial_clause_prev[9][33] & 1'b1;
			partial_clause[9][34] 	= partial_clause_prev[9][34] & 1'b1;
			partial_clause[9][35] 	= partial_clause_prev[9][35] & 1'b1;
			partial_clause[9][36] 	= partial_clause_prev[9][36] & 1'b1;
			partial_clause[9][37] 	= partial_clause_prev[9][37] & 1'b1;
			partial_clause[9][38] 	= partial_clause_prev[9][38] & 1'b1;
			partial_clause[9][39] 	= partial_clause_prev[9][39] & ~x[5];
			partial_clause[9][40] 	= partial_clause_prev[9][40] & 1'b1;
			partial_clause[9][41] 	= partial_clause_prev[9][41] & 1'b1;
			partial_clause[9][42] 	= partial_clause_prev[9][42] & 1'b1;
			partial_clause[9][43] 	= partial_clause_prev[9][43] & 1'b1;
			partial_clause[9][44] 	= partial_clause_prev[9][44] & 1'b1;
			partial_clause[9][45] 	= partial_clause_prev[9][45] & 1'b1;
			partial_clause[9][46] 	= partial_clause_prev[9][46] & 1'b1;
			partial_clause[9][47] 	= partial_clause_prev[9][47] & 1'b1;
			partial_clause[9][48] 	= partial_clause_prev[9][48] & 1'b1;
			partial_clause[9][49] 	= partial_clause_prev[9][49] & 1'b1;
			partial_clause[9][50] 	= partial_clause_prev[9][50] & 1'b1;
			partial_clause[9][51] 	= partial_clause_prev[9][51] & 1'b1;
			partial_clause[9][52] 	= partial_clause_prev[9][52] & 1'b1;
			partial_clause[9][53] 	= partial_clause_prev[9][53] & ~x[13];
			partial_clause[9][54] 	= partial_clause_prev[9][54] & 1'b1;
			partial_clause[9][55] 	= partial_clause_prev[9][55] & 1'b1;
			partial_clause[9][56] 	= partial_clause_prev[9][56] & ~x[5];
			partial_clause[9][57] 	= partial_clause_prev[9][57] & 1'b1;
			partial_clause[9][58] 	= partial_clause_prev[9][58] & 1'b1;
			partial_clause[9][59] 	= partial_clause_prev[9][59] & 1'b1;
			partial_clause[9][60] 	= partial_clause_prev[9][60] & 1'b1;
			partial_clause[9][61] 	= partial_clause_prev[9][61] & 1'b1;
			partial_clause[9][62] 	= partial_clause_prev[9][62] & 1'b1;
			partial_clause[9][63] 	= partial_clause_prev[9][63] & 1'b1;
			partial_clause[9][64] 	= partial_clause_prev[9][64] & 1'b1;
			partial_clause[9][65] 	= partial_clause_prev[9][65] & 1'b1;
			partial_clause[9][66] 	= partial_clause_prev[9][66] & 1'b1;
			partial_clause[9][67] 	= partial_clause_prev[9][67] & 1'b1;
			partial_clause[9][68] 	= partial_clause_prev[9][68] & 1'b1;
			partial_clause[9][69] 	= partial_clause_prev[9][69] & 1'b1;
			partial_clause[9][70] 	= partial_clause_prev[9][70] & 1'b1;
			partial_clause[9][71] 	= partial_clause_prev[9][71] & 1'b1;
			partial_clause[9][72] 	= partial_clause_prev[9][72] & ~x[7];
			partial_clause[9][73] 	= partial_clause_prev[9][73] & 1'b1;
			partial_clause[9][74] 	= partial_clause_prev[9][74] & 1'b1;
			partial_clause[9][75] 	= partial_clause_prev[9][75] & ~x[9];
			partial_clause[9][76] 	= partial_clause_prev[9][76] & 1'b1;
			partial_clause[9][77] 	= partial_clause_prev[9][77] & 1'b1;
			partial_clause[9][78] 	= partial_clause_prev[9][78] & 1'b1;
			partial_clause[9][79] 	= partial_clause_prev[9][79] & 1'b1;
			partial_clause[9][80] 	= partial_clause_prev[9][80] & 1'b1;
			partial_clause[9][81] 	= partial_clause_prev[9][81] & 1'b1;
			partial_clause[9][82] 	= partial_clause_prev[9][82] & 1'b1;
			partial_clause[9][83] 	= partial_clause_prev[9][83] & ~x[2];
			partial_clause[9][84] 	= partial_clause_prev[9][84] & 1'b1;
			partial_clause[9][85] 	= partial_clause_prev[9][85] & 1'b1;
			partial_clause[9][86] 	= partial_clause_prev[9][86] & 1'b1;
			partial_clause[9][87] 	= partial_clause_prev[9][87] & 1'b1;
			partial_clause[9][88] 	= partial_clause_prev[9][88] & 1'b1;
			partial_clause[9][89] 	= partial_clause_prev[9][89] & 1'b1;
			partial_clause[9][90] 	= partial_clause_prev[9][90] & 1'b1;
			partial_clause[9][91] 	= partial_clause_prev[9][91] & 1'b1;
			partial_clause[9][92] 	= partial_clause_prev[9][92] & 1'b1;
			partial_clause[9][93] 	= partial_clause_prev[9][93] & 1'b1;
			partial_clause[9][94] 	= partial_clause_prev[9][94] & 1'b1;
			partial_clause[9][95] 	= partial_clause_prev[9][95] & 1'b1;
			partial_clause[9][96] 	= partial_clause_prev[9][96] & 1'b1;
			partial_clause[9][97] 	= partial_clause_prev[9][97] & 1'b1;
			partial_clause[9][98] 	= partial_clause_prev[9][98] & 1'b1;
			partial_clause[9][99] 	= partial_clause_prev[9][99] & 1'b1;
		end
	end
endmodule


