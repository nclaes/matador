module HCB_0 (x, partial_clause, clk, valid);
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= ~x[2] & ~x[6] & ~x[9] & ~x[13] & ~x[14] & ~x[17] & ~x[23] & ~x[27] & ~x[28] & ~x[30] & ~x[33] & ~x[34] & ~x[39] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[45] & ~x[47] & ~x[50] & ~x[57] & ~x[59] & ~x[63];
			partial_clause[1] 	= ~x[8] & ~x[20] & ~x[22] & ~x[27] & ~x[31] & ~x[43] & ~x[61] & ~x[63];
			partial_clause[2] 	= ~x[1] & ~x[7] & ~x[10] & ~x[27];
			partial_clause[3] 	= ~x[9] & ~x[13] & ~x[32] & ~x[33] & ~x[37] & ~x[42] & ~x[58];
			partial_clause[4] 	= ~x[1] & ~x[5] & ~x[19] & ~x[24] & ~x[28] & ~x[33] & ~x[49] & ~x[52] & ~x[54];
			partial_clause[5] 	= ~x[1] & ~x[3] & ~x[4] & ~x[6] & ~x[10] & ~x[17] & ~x[24] & ~x[28] & ~x[33] & ~x[37] & ~x[47] & ~x[54] & ~x[58];
			partial_clause[6] 	= ~x[1] & ~x[14] & ~x[21] & ~x[42] & ~x[61];
			partial_clause[7] 	= ~x[0] & ~x[3] & ~x[9] & ~x[11] & ~x[13] & ~x[15] & ~x[25] & ~x[26] & ~x[47];
			partial_clause[8] 	= ~x[1] & ~x[10] & ~x[24] & ~x[33] & ~x[34] & ~x[35] & ~x[39] & ~x[50] & ~x[51] & ~x[57] & ~x[61];
			partial_clause[9] 	= ~x[2] & ~x[6] & ~x[18] & ~x[22] & ~x[23] & ~x[27] & ~x[29] & ~x[32] & ~x[33] & ~x[34] & ~x[37] & ~x[43] & ~x[46] & ~x[47] & ~x[51] & ~x[52] & ~x[55] & ~x[56] & ~x[61];
			partial_clause[10] 	= ~x[2] & ~x[5] & ~x[10] & ~x[14] & ~x[27] & ~x[28] & ~x[29] & ~x[31] & ~x[32] & ~x[35] & ~x[41] & ~x[49] & ~x[54] & ~x[58] & ~x[59] & ~x[61];
			partial_clause[11] 	= ~x[17] & ~x[18] & ~x[22] & ~x[23] & ~x[28] & ~x[35] & ~x[40] & ~x[41] & ~x[43] & ~x[50] & ~x[52] & ~x[60] & ~x[61];
			partial_clause[12] 	= ~x[1] & ~x[3] & ~x[7] & ~x[13] & ~x[26] & ~x[33] & ~x[36] & ~x[38] & ~x[39] & ~x[40] & ~x[46] & ~x[49] & ~x[50] & ~x[56] & ~x[62];
			partial_clause[13] 	= ~x[0] & ~x[4] & ~x[6] & ~x[10] & ~x[17] & ~x[33] & ~x[34] & ~x[37] & ~x[41] & ~x[52] & ~x[54] & ~x[63];
			partial_clause[14] 	= ~x[20];
			partial_clause[15] 	= 1'b1;
			partial_clause[16] 	= ~x[12] & ~x[26] & ~x[31] & ~x[37] & ~x[56] & ~x[58];
			partial_clause[17] 	= 1'b1;
			partial_clause[18] 	= ~x[15] & ~x[23] & ~x[29] & ~x[36] & ~x[45] & ~x[62];
			partial_clause[19] 	= ~x[9] & ~x[16] & ~x[24] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & ~x[30] & ~x[34] & ~x[50] & ~x[54] & ~x[58] & ~x[59] & ~x[61];
			partial_clause[20] 	= ~x[3] & ~x[23] & ~x[41];
			partial_clause[21] 	= ~x[5] & ~x[40] & ~x[57] & ~x[60];
			partial_clause[22] 	= ~x[2] & ~x[14] & ~x[22];
			partial_clause[23] 	= ~x[3] & ~x[4] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[12] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[23] & ~x[24] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[35] & ~x[36] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[45] & ~x[46] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[59] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[24] 	= ~x[2] & ~x[3] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[11] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[19] & ~x[22] & ~x[25] & ~x[26] & ~x[27] & ~x[30] & ~x[32] & ~x[35] & ~x[37] & ~x[38] & ~x[40] & ~x[43] & ~x[44] & ~x[45] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[53] & ~x[54] & ~x[57] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[25] 	= ~x[0] & ~x[5] & ~x[8] & ~x[9] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[19] & ~x[22] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & ~x[30] & ~x[32] & ~x[45] & ~x[46] & ~x[48] & ~x[51] & ~x[54] & ~x[56] & ~x[57] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[26] 	= 1'b1;
			partial_clause[27] 	= ~x[10] & ~x[11] & ~x[16] & ~x[28] & ~x[34] & ~x[45] & ~x[49] & ~x[61];
			partial_clause[28] 	= ~x[4] & ~x[14] & ~x[16] & ~x[25] & ~x[35] & ~x[36] & ~x[41] & ~x[55];
			partial_clause[29] 	= ~x[15] & ~x[31] & ~x[33] & ~x[38] & ~x[40] & ~x[62];
			partial_clause[30] 	= ~x[13] & ~x[32] & ~x[34] & ~x[39] & ~x[46] & ~x[47] & ~x[61];
			partial_clause[31] 	= ~x[4] & ~x[22] & ~x[34] & ~x[58] & ~x[60];
			partial_clause[32] 	= ~x[0] & ~x[13] & ~x[17] & ~x[29] & ~x[38];
			partial_clause[33] 	= 1'b1;
			partial_clause[34] 	= ~x[2] & ~x[3] & ~x[6] & ~x[8] & ~x[11] & ~x[14] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[27] & ~x[30] & ~x[36] & ~x[39] & ~x[40] & ~x[41] & ~x[42] & ~x[46] & ~x[53] & ~x[56] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[35] 	= ~x[35] & ~x[53];
			partial_clause[36] 	= ~x[0] & ~x[4] & ~x[5] & ~x[11] & ~x[22] & ~x[27] & ~x[41] & ~x[52] & ~x[53] & ~x[54];
			partial_clause[37] 	= ~x[8] & ~x[13] & ~x[24] & ~x[32] & ~x[42] & ~x[51] & ~x[56];
			partial_clause[38] 	= ~x[7] & ~x[20] & ~x[24] & ~x[27] & ~x[28] & ~x[33] & ~x[40] & ~x[49] & ~x[50] & ~x[54] & ~x[55] & ~x[62];
			partial_clause[39] 	= ~x[0] & ~x[5] & ~x[8] & ~x[42];
			partial_clause[40] 	= ~x[6] & ~x[17] & ~x[20] & ~x[45] & ~x[57];
			partial_clause[41] 	= 1'b1;
			partial_clause[42] 	= ~x[14] & ~x[16] & ~x[22] & ~x[24] & ~x[37] & ~x[42] & ~x[61];
			partial_clause[43] 	= ~x[7] & ~x[11] & ~x[13] & ~x[33] & ~x[47] & ~x[61];
			partial_clause[44] 	= 1'b1;
			partial_clause[45] 	= ~x[48];
			partial_clause[46] 	= ~x[0] & ~x[3] & ~x[5] & ~x[10] & ~x[12] & ~x[18] & ~x[24] & ~x[30] & ~x[35] & ~x[36] & ~x[38] & ~x[41] & ~x[44] & ~x[45] & ~x[48] & ~x[49] & ~x[52] & ~x[53] & ~x[54] & ~x[57] & ~x[61];
			partial_clause[47] 	= ~x[16] & ~x[23] & ~x[34] & ~x[46] & ~x[54] & ~x[55];
			partial_clause[48] 	= 1'b1;
			partial_clause[49] 	= 1'b1;
			partial_clause[50] 	= ~x[1] & ~x[7] & ~x[16] & ~x[25] & ~x[30] & ~x[36] & ~x[39] & ~x[48] & ~x[54];
			partial_clause[51] 	= 1'b1;
			partial_clause[52] 	= 1'b1;
			partial_clause[53] 	= 1'b1;
			partial_clause[54] 	= ~x[30];
			partial_clause[55] 	= ~x[5];
			partial_clause[56] 	= 1'b1;
			partial_clause[57] 	= ~x[1] & ~x[11] & ~x[27] & ~x[29] & ~x[31] & ~x[39] & ~x[51] & ~x[54] & ~x[58] & ~x[61];
			partial_clause[58] 	= ~x[8] & ~x[15] & ~x[32] & ~x[53] & ~x[56] & ~x[57];
			partial_clause[59] 	= ~x[8] & ~x[9] & ~x[15] & ~x[23] & ~x[29] & ~x[31] & ~x[41] & ~x[48] & ~x[57] & ~x[60] & ~x[61];
			partial_clause[60] 	= 1'b1;
			partial_clause[61] 	= ~x[62];
			partial_clause[62] 	= ~x[9] & ~x[14] & ~x[15] & ~x[20] & ~x[21] & ~x[25] & ~x[34] & ~x[40] & ~x[48] & ~x[52];
			partial_clause[63] 	= ~x[3] & ~x[36];
			partial_clause[64] 	= 1'b1;
			partial_clause[65] 	= 1'b1;
			partial_clause[66] 	= 1'b1;
			partial_clause[67] 	= 1'b1;
			partial_clause[68] 	= ~x[10] & ~x[20] & ~x[26] & ~x[27] & ~x[39] & ~x[40];
			partial_clause[69] 	= ~x[5] & ~x[34] & ~x[43] & ~x[55];
			partial_clause[70] 	= ~x[4] & ~x[9] & ~x[21] & ~x[23] & ~x[27] & ~x[31] & ~x[53] & ~x[60];
			partial_clause[71] 	= ~x[46];
			partial_clause[72] 	= 1'b1;
			partial_clause[73] 	= ~x[38];
			partial_clause[74] 	= ~x[5] & ~x[11] & ~x[27] & ~x[32] & ~x[35] & ~x[41] & ~x[43] & ~x[47];
			partial_clause[75] 	= ~x[3] & ~x[39] & ~x[42] & ~x[43];
			partial_clause[76] 	= ~x[3] & ~x[12] & ~x[15] & ~x[20] & ~x[22] & ~x[24] & ~x[27] & ~x[38] & ~x[43] & ~x[44] & ~x[45] & ~x[53] & ~x[54] & ~x[56] & ~x[58] & ~x[59];
			partial_clause[77] 	= ~x[9] & ~x[11] & ~x[14] & ~x[44];
			partial_clause[78] 	= ~x[16];
			partial_clause[79] 	= ~x[0] & ~x[10] & ~x[15] & ~x[24] & ~x[59];
			partial_clause[80] 	= 1'b1;
			partial_clause[81] 	= ~x[1];
			partial_clause[82] 	= 1'b1;
			partial_clause[83] 	= 1'b1;
			partial_clause[84] 	= ~x[1] & ~x[13] & ~x[36];
			partial_clause[85] 	= ~x[0] & ~x[3] & ~x[5] & ~x[7] & ~x[17] & ~x[26] & ~x[31] & ~x[48] & ~x[49] & ~x[56];
			partial_clause[86] 	= ~x[3] & ~x[7] & ~x[30] & ~x[32] & ~x[36] & ~x[50] & ~x[58];
			partial_clause[87] 	= ~x[10] & ~x[13] & ~x[18] & ~x[55] & ~x[63];
			partial_clause[88] 	= ~x[7] & ~x[8] & ~x[12] & ~x[17] & ~x[18] & ~x[19] & ~x[21] & ~x[24] & ~x[28] & ~x[35] & ~x[37] & ~x[63];
			partial_clause[89] 	= ~x[3] & ~x[5] & ~x[16] & ~x[20] & ~x[49];
			partial_clause[90] 	= 1'b1;
			partial_clause[91] 	= ~x[4] & ~x[30];
			partial_clause[92] 	= ~x[48];
			partial_clause[93] 	= ~x[1] & ~x[2] & ~x[4] & ~x[5] & ~x[11] & ~x[15] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[34] & ~x[35] & ~x[38] & ~x[39] & ~x[44] & ~x[47] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[59] & ~x[62] & ~x[63];
			partial_clause[94] 	= 1'b1;
			partial_clause[95] 	= ~x[1] & ~x[3] & ~x[4] & ~x[8] & ~x[11] & ~x[13] & ~x[29] & ~x[32] & ~x[36] & ~x[37] & ~x[44] & ~x[49] & ~x[50];
			partial_clause[96] 	= ~x[4];
			partial_clause[97] 	= ~x[4] & ~x[8] & ~x[16] & ~x[20] & ~x[26] & ~x[27] & ~x[29] & ~x[34] & ~x[41] & ~x[43] & ~x[45] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[57] & ~x[58] & ~x[62] & ~x[63];
			partial_clause[98] 	= ~x[3] & ~x[5] & ~x[7] & ~x[9] & ~x[12] & ~x[24] & ~x[31] & ~x[41] & ~x[51] & ~x[57] & ~x[58] & ~x[59] & ~x[62];
			partial_clause[99] 	= ~x[0] & ~x[1] & ~x[2] & ~x[4] & ~x[9] & ~x[10] & ~x[13] & ~x[14] & ~x[15] & ~x[18] & ~x[20] & ~x[22] & ~x[27] & ~x[30] & ~x[33] & ~x[35] & ~x[39] & ~x[41] & ~x[43] & ~x[44] & ~x[47] & ~x[50] & ~x[51] & ~x[53] & ~x[56] & ~x[57] & ~x[58] & ~x[59] & ~x[61] & ~x[63];
			partial_clause[100] 	= ~x[48] & ~x[51] & ~x[52];
			partial_clause[101] 	= ~x[9] & ~x[39];
			partial_clause[102] 	= ~x[7] & ~x[13];
			partial_clause[103] 	= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[10] & ~x[13] & ~x[15] & ~x[16] & ~x[19] & ~x[22] & ~x[30] & ~x[33] & ~x[34] & ~x[35] & ~x[37] & ~x[41] & ~x[47] & ~x[50] & ~x[51] & ~x[55] & ~x[57] & ~x[62];
			partial_clause[104] 	= ~x[1] & ~x[4] & ~x[19] & ~x[41] & ~x[50];
			partial_clause[105] 	= ~x[0] & ~x[3] & ~x[4] & ~x[7] & ~x[13] & ~x[14] & ~x[21] & ~x[24] & ~x[26] & ~x[27] & ~x[30] & ~x[32] & ~x[33] & ~x[37] & ~x[45] & ~x[48] & ~x[51] & ~x[59] & ~x[60] & ~x[62];
			partial_clause[106] 	= ~x[4] & ~x[15] & ~x[25] & ~x[31] & ~x[41] & ~x[56];
			partial_clause[107] 	= ~x[2] & ~x[6] & ~x[7] & ~x[15] & ~x[17] & ~x[20] & ~x[22] & ~x[27] & ~x[32] & ~x[34] & ~x[37] & ~x[42] & ~x[48] & ~x[49] & ~x[50];
			partial_clause[108] 	= ~x[4] & ~x[9] & ~x[14] & ~x[15] & ~x[16] & ~x[19] & ~x[24] & ~x[29] & ~x[33] & ~x[34] & ~x[38] & ~x[39] & ~x[42] & ~x[48] & ~x[54] & ~x[61];
			partial_clause[109] 	= 1'b1;
			partial_clause[110] 	= ~x[19];
			partial_clause[111] 	= 1'b1;
			partial_clause[112] 	= ~x[3] & ~x[10] & ~x[27] & ~x[49];
			partial_clause[113] 	= ~x[12] & ~x[39] & ~x[43] & ~x[47] & ~x[59];
			partial_clause[114] 	= 1'b1;
			partial_clause[115] 	= ~x[1] & ~x[5] & ~x[10] & ~x[11] & ~x[14] & ~x[18] & ~x[19] & ~x[21] & ~x[23] & ~x[24] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[44] & ~x[46] & ~x[49] & ~x[51] & ~x[53] & ~x[55] & ~x[60];
			partial_clause[116] 	= ~x[5] & ~x[19] & ~x[22] & ~x[28] & ~x[37] & ~x[42] & ~x[45];
			partial_clause[117] 	= 1'b1;
			partial_clause[118] 	= ~x[6] & ~x[7] & ~x[12] & ~x[25] & ~x[26] & ~x[34] & ~x[35] & ~x[41] & ~x[42] & ~x[44] & ~x[56] & ~x[61];
			partial_clause[119] 	= ~x[2] & ~x[12] & ~x[15] & ~x[17] & ~x[20] & ~x[21] & ~x[23] & ~x[25] & ~x[26] & ~x[27] & ~x[32] & ~x[33] & ~x[34] & ~x[35] & ~x[41] & ~x[44] & ~x[54] & ~x[61] & ~x[63];
			partial_clause[120] 	= ~x[1] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[15] & ~x[16] & ~x[17] & ~x[19] & ~x[21] & ~x[22] & ~x[23] & ~x[25] & ~x[26] & ~x[32] & ~x[35] & ~x[38] & ~x[39] & ~x[40] & ~x[41] & ~x[45] & ~x[46] & ~x[48] & ~x[50] & ~x[51] & ~x[52] & ~x[54] & ~x[55] & ~x[57] & ~x[58] & ~x[59] & ~x[62];
			partial_clause[121] 	= ~x[6] & ~x[11] & ~x[14] & ~x[22] & ~x[24] & ~x[25] & ~x[29] & ~x[30] & ~x[35] & ~x[47] & ~x[50] & ~x[60];
			partial_clause[122] 	= ~x[11] & ~x[29] & ~x[41] & ~x[48] & ~x[50];
			partial_clause[123] 	= ~x[0] & ~x[8] & ~x[10] & ~x[12] & ~x[17] & ~x[19] & ~x[20] & ~x[22] & ~x[23] & ~x[28] & ~x[31] & ~x[32] & ~x[34] & ~x[41] & ~x[42] & ~x[45] & ~x[53] & ~x[55] & ~x[58];
			partial_clause[124] 	= 1'b1;
			partial_clause[125] 	= ~x[4] & ~x[24] & ~x[31] & ~x[38] & ~x[43] & ~x[48] & ~x[61];
			partial_clause[126] 	= ~x[14] & ~x[15] & ~x[50];
			partial_clause[127] 	= ~x[1] & ~x[8] & ~x[10] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[23] & ~x[25] & ~x[26] & ~x[27] & ~x[30] & ~x[31] & ~x[32] & ~x[34] & ~x[35] & ~x[38] & ~x[39] & ~x[40] & ~x[43] & ~x[44] & ~x[46] & ~x[49] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[56] & ~x[59] & ~x[63];
			partial_clause[128] 	= ~x[4] & ~x[9] & ~x[15] & ~x[31];
			partial_clause[129] 	= ~x[4] & ~x[9] & ~x[11] & ~x[12] & ~x[17] & ~x[18] & ~x[24] & ~x[26] & ~x[27] & ~x[32] & ~x[43] & ~x[44] & ~x[46] & ~x[51] & ~x[52] & ~x[57] & ~x[59] & ~x[60];
			partial_clause[130] 	= ~x[9] & ~x[14] & ~x[23] & ~x[26] & ~x[28] & ~x[33] & ~x[36] & ~x[43] & ~x[52] & ~x[58] & ~x[63];
			partial_clause[131] 	= ~x[60] & ~x[61];
			partial_clause[132] 	= ~x[24] & ~x[32] & ~x[46];
			partial_clause[133] 	= ~x[2] & ~x[61];
			partial_clause[134] 	= ~x[1] & ~x[5] & ~x[6] & ~x[13] & ~x[17] & ~x[21] & ~x[24] & ~x[32] & ~x[37] & ~x[39] & ~x[42] & ~x[43] & ~x[48] & ~x[50] & ~x[54] & ~x[56] & ~x[57] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[135] 	= ~x[12] & ~x[24] & ~x[31] & ~x[41] & ~x[45] & ~x[57];
			partial_clause[136] 	= ~x[1] & ~x[3] & ~x[8] & ~x[9] & ~x[11] & ~x[14] & ~x[23] & ~x[25] & ~x[26] & ~x[31] & ~x[43] & ~x[50] & ~x[51] & ~x[55] & ~x[57] & ~x[63];
			partial_clause[137] 	= 1'b1;
			partial_clause[138] 	= 1'b1;
			partial_clause[139] 	= ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[23] & ~x[25] & ~x[27] & ~x[30] & ~x[34] & ~x[43] & ~x[48] & ~x[51] & ~x[53] & ~x[60] & ~x[63];
			partial_clause[140] 	= ~x[2] & ~x[5] & ~x[7] & ~x[18] & ~x[19] & ~x[20] & ~x[24] & ~x[25] & ~x[30] & ~x[31] & ~x[32] & ~x[34] & ~x[36] & ~x[37] & ~x[39] & ~x[44] & ~x[50] & ~x[56] & ~x[58];
			partial_clause[141] 	= ~x[61];
			partial_clause[142] 	= ~x[3] & ~x[4] & ~x[12] & ~x[13] & ~x[24] & ~x[33] & ~x[39] & ~x[40] & ~x[41] & ~x[42] & ~x[49] & ~x[50] & ~x[55] & ~x[56] & ~x[59];
			partial_clause[143] 	= 1'b1;
			partial_clause[144] 	= ~x[2] & ~x[15] & ~x[22] & ~x[26] & ~x[27] & ~x[37] & ~x[39] & ~x[44] & ~x[46] & ~x[47] & ~x[55];
			partial_clause[145] 	= 1'b1;
			partial_clause[146] 	= ~x[5] & ~x[11] & ~x[16] & ~x[21] & ~x[53] & ~x[63];
			partial_clause[147] 	= ~x[20] & ~x[22] & ~x[23] & ~x[24] & ~x[31] & ~x[32] & ~x[43] & ~x[50] & ~x[56] & ~x[58] & ~x[59] & ~x[63];
			partial_clause[148] 	= ~x[3] & ~x[15] & ~x[18] & ~x[19] & ~x[42] & ~x[50] & ~x[58];
			partial_clause[149] 	= ~x[21] & ~x[26] & ~x[48];
			partial_clause[150] 	= ~x[3] & ~x[4] & ~x[12] & ~x[18] & ~x[41] & ~x[49] & ~x[52] & ~x[54] & ~x[55];
			partial_clause[151] 	= ~x[2];
			partial_clause[152] 	= ~x[11] & ~x[13] & ~x[15] & ~x[16] & ~x[27] & ~x[44] & ~x[53];
			partial_clause[153] 	= ~x[10] & ~x[11] & ~x[15] & ~x[29] & ~x[32] & ~x[38] & ~x[47] & ~x[48] & ~x[52] & ~x[62];
			partial_clause[154] 	= ~x[40] & ~x[56];
			partial_clause[155] 	= 1'b1;
			partial_clause[156] 	= ~x[21];
			partial_clause[157] 	= 1'b1;
			partial_clause[158] 	= ~x[0] & ~x[4] & ~x[6] & ~x[9] & ~x[11] & ~x[12] & ~x[16] & ~x[18] & ~x[20] & ~x[24] & ~x[25] & ~x[27] & ~x[28] & ~x[30] & ~x[31] & ~x[35] & ~x[36] & ~x[37] & ~x[43] & ~x[47] & ~x[49] & ~x[51] & ~x[52] & ~x[53] & ~x[54] & ~x[58] & ~x[59] & ~x[62];
			partial_clause[159] 	= ~x[9] & ~x[16] & ~x[18] & ~x[24] & ~x[27] & ~x[31] & ~x[38] & ~x[39] & ~x[41] & ~x[42] & ~x[46] & ~x[56];
			partial_clause[160] 	= ~x[0] & ~x[8] & ~x[22] & ~x[42] & ~x[57] & ~x[63];
			partial_clause[161] 	= ~x[3] & ~x[16] & ~x[25] & ~x[28] & ~x[32] & ~x[33] & ~x[39] & ~x[42] & ~x[45] & ~x[49] & ~x[51] & ~x[55];
			partial_clause[162] 	= ~x[2] & ~x[6] & ~x[10] & ~x[32] & ~x[42];
			partial_clause[163] 	= 1'b1;
			partial_clause[164] 	= ~x[1] & ~x[16] & ~x[18] & ~x[54] & ~x[61];
			partial_clause[165] 	= ~x[1] & ~x[8] & ~x[14] & ~x[20] & ~x[21] & ~x[22] & ~x[25] & ~x[30] & ~x[48] & ~x[51] & ~x[52] & ~x[58] & ~x[60];
			partial_clause[166] 	= ~x[0] & ~x[2] & ~x[9] & ~x[17] & ~x[23] & ~x[24] & ~x[26] & ~x[34] & ~x[38] & ~x[43] & ~x[46] & ~x[51] & ~x[56] & ~x[60];
			partial_clause[167] 	= 1'b1;
			partial_clause[168] 	= ~x[16] & ~x[46];
			partial_clause[169] 	= ~x[0] & ~x[7] & ~x[18] & ~x[37] & ~x[51];
			partial_clause[170] 	= 1'b1;
			partial_clause[171] 	= ~x[2] & ~x[4] & ~x[5] & ~x[19] & ~x[26] & ~x[39] & ~x[41] & ~x[44] & ~x[49] & ~x[53] & ~x[62];
			partial_clause[172] 	= 1'b1;
			partial_clause[173] 	= ~x[9] & ~x[10] & ~x[14] & ~x[16] & ~x[24] & ~x[41] & ~x[43] & ~x[56] & ~x[60] & ~x[61];
			partial_clause[174] 	= ~x[48] & ~x[60];
			partial_clause[175] 	= 1'b1;
			partial_clause[176] 	= ~x[1] & ~x[18] & ~x[35] & ~x[43];
			partial_clause[177] 	= ~x[10] & ~x[33] & ~x[54];
			partial_clause[178] 	= ~x[12] & ~x[19] & ~x[48] & ~x[55] & ~x[61];
			partial_clause[179] 	= ~x[29] & ~x[60];
			partial_clause[180] 	= ~x[34] & ~x[52] & ~x[58];
			partial_clause[181] 	= 1'b1;
			partial_clause[182] 	= 1'b1;
			partial_clause[183] 	= ~x[0] & ~x[7] & ~x[11] & ~x[14] & ~x[15] & ~x[18] & ~x[21] & ~x[22] & ~x[24] & ~x[31] & ~x[33] & ~x[34] & ~x[38] & ~x[47] & ~x[58] & ~x[59] & ~x[63];
			partial_clause[184] 	= ~x[0] & ~x[7] & ~x[11] & ~x[17] & ~x[21] & ~x[23] & ~x[25] & ~x[26] & ~x[33] & ~x[49] & ~x[51] & ~x[53] & ~x[55] & ~x[58] & ~x[60] & ~x[62];
			partial_clause[185] 	= ~x[3] & ~x[4] & ~x[6] & ~x[32] & ~x[56] & ~x[63];
			partial_clause[186] 	= ~x[0] & ~x[3] & ~x[15] & ~x[16] & ~x[18] & ~x[19] & ~x[28] & ~x[33] & ~x[34] & ~x[37] & ~x[50] & ~x[51] & ~x[53] & ~x[59] & ~x[60];
			partial_clause[187] 	= ~x[4] & ~x[5] & ~x[12] & ~x[16] & ~x[23] & ~x[28] & ~x[29] & ~x[30] & ~x[35] & ~x[48] & ~x[53] & ~x[54] & ~x[58];
			partial_clause[188] 	= ~x[16];
			partial_clause[189] 	= 1'b1;
			partial_clause[190] 	= ~x[10] & ~x[26] & ~x[32] & ~x[37] & ~x[39] & ~x[44] & ~x[59];
			partial_clause[191] 	= ~x[27];
			partial_clause[192] 	= ~x[32] & ~x[33];
			partial_clause[193] 	= ~x[2] & ~x[16] & ~x[30] & ~x[40];
			partial_clause[194] 	= ~x[5] & ~x[9];
			partial_clause[195] 	= ~x[5] & ~x[7] & ~x[10] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[17] & ~x[24] & ~x[25] & ~x[26] & ~x[35] & ~x[40] & ~x[44] & ~x[45] & ~x[46] & ~x[50] & ~x[53] & ~x[55] & ~x[62] & ~x[63];
			partial_clause[196] 	= ~x[47] & ~x[49];
			partial_clause[197] 	= ~x[5] & ~x[11] & ~x[12] & ~x[13] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[29] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[34] & ~x[38] & ~x[46] & ~x[47] & ~x[51];
			partial_clause[198] 	= ~x[49];
			partial_clause[199] 	= 1'b1;
			partial_clause[200] 	= ~x[9] & ~x[14] & ~x[18] & ~x[28] & ~x[63];
			partial_clause[201] 	= ~x[4] & ~x[8] & ~x[18] & ~x[32] & ~x[34] & ~x[46] & ~x[51] & ~x[54] & ~x[62];
			partial_clause[202] 	= ~x[1] & ~x[2] & ~x[10] & ~x[15] & ~x[19] & ~x[22] & ~x[23] & ~x[27] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[34] & ~x[40] & ~x[41] & ~x[49] & ~x[52] & ~x[53] & ~x[56] & ~x[57] & ~x[58];
			partial_clause[203] 	= ~x[11];
			partial_clause[204] 	= ~x[9] & ~x[10] & ~x[18] & ~x[21] & ~x[25] & ~x[26] & ~x[27] & ~x[28] & ~x[31] & ~x[36] & ~x[40] & ~x[43] & ~x[50] & ~x[51] & ~x[54] & ~x[57] & ~x[61];
			partial_clause[205] 	= 1'b1;
			partial_clause[206] 	= ~x[2] & ~x[4] & ~x[12] & ~x[13] & ~x[18] & ~x[32] & ~x[35] & ~x[40] & ~x[43] & ~x[44] & ~x[46] & ~x[49] & ~x[54] & ~x[55] & ~x[59] & ~x[60] & ~x[63];
			partial_clause[207] 	= ~x[39] & ~x[55] & ~x[56];
			partial_clause[208] 	= ~x[10] & ~x[20] & ~x[22] & ~x[30] & ~x[33] & ~x[48];
			partial_clause[209] 	= ~x[43];
			partial_clause[210] 	= ~x[2] & ~x[3] & ~x[18] & ~x[22] & ~x[35] & ~x[61];
			partial_clause[211] 	= 1'b1;
			partial_clause[212] 	= ~x[15] & ~x[18] & ~x[25];
			partial_clause[213] 	= 1'b1;
			partial_clause[214] 	= 1'b1;
			partial_clause[215] 	= 1'b1;
			partial_clause[216] 	= ~x[30] & ~x[35];
			partial_clause[217] 	= ~x[8] & ~x[21] & ~x[26] & ~x[27] & ~x[38] & ~x[40] & ~x[44];
			partial_clause[218] 	= ~x[55];
			partial_clause[219] 	= ~x[15] & ~x[24] & ~x[28] & ~x[43] & ~x[48] & ~x[50];
			partial_clause[220] 	= ~x[1] & ~x[3] & ~x[4] & ~x[5] & ~x[7] & ~x[8] & ~x[11] & ~x[13] & ~x[14] & ~x[16] & ~x[20] & ~x[21] & ~x[25] & ~x[30] & ~x[31] & ~x[36] & ~x[42] & ~x[49] & ~x[50] & ~x[52] & ~x[55] & ~x[56] & ~x[57] & ~x[59];
			partial_clause[221] 	= 1'b1;
			partial_clause[222] 	= 1'b1;
			partial_clause[223] 	= ~x[7] & ~x[26] & ~x[34] & ~x[39] & ~x[42] & ~x[43];
			partial_clause[224] 	= ~x[3] & ~x[11] & ~x[16] & ~x[19] & ~x[20] & ~x[24] & ~x[25] & ~x[44] & ~x[57] & ~x[60];
			partial_clause[225] 	= ~x[40] & ~x[59];
			partial_clause[226] 	= ~x[1] & ~x[3] & ~x[6] & ~x[11] & ~x[13] & ~x[16] & ~x[17] & ~x[19] & ~x[21] & ~x[23] & ~x[25] & ~x[28] & ~x[30] & ~x[33] & ~x[40] & ~x[45] & ~x[46] & ~x[48] & ~x[50] & ~x[51] & ~x[57] & ~x[62];
			partial_clause[227] 	= ~x[13] & ~x[49] & ~x[55];
			partial_clause[228] 	= ~x[17] & ~x[21] & ~x[32] & ~x[34] & ~x[43] & ~x[46] & ~x[49] & ~x[62] & ~x[63];
			partial_clause[229] 	= ~x[2] & ~x[25] & ~x[34] & ~x[36] & ~x[37] & ~x[38] & ~x[39] & ~x[41] & ~x[45] & ~x[46] & ~x[52] & ~x[53] & ~x[57] & ~x[60];
			partial_clause[230] 	= ~x[1] & ~x[2] & ~x[5] & ~x[6] & ~x[8] & ~x[15] & ~x[19] & ~x[27] & ~x[28] & ~x[30] & ~x[31] & ~x[38] & ~x[40] & ~x[43] & ~x[45] & ~x[47] & ~x[50] & ~x[52] & ~x[56] & ~x[58] & ~x[62];
			partial_clause[231] 	= ~x[1] & ~x[5] & ~x[12] & ~x[21] & ~x[28] & ~x[47] & ~x[48] & ~x[53];
			partial_clause[232] 	= 1'b1;
			partial_clause[233] 	= ~x[2] & ~x[21] & ~x[28] & ~x[40] & ~x[42] & ~x[56] & ~x[60];
			partial_clause[234] 	= ~x[29] & ~x[34];
			partial_clause[235] 	= 1'b1;
			partial_clause[236] 	= 1'b1;
			partial_clause[237] 	= ~x[27];
			partial_clause[238] 	= ~x[17] & ~x[25];
			partial_clause[239] 	= ~x[21] & ~x[26] & ~x[57];
			partial_clause[240] 	= ~x[4] & ~x[6] & ~x[17] & ~x[20] & ~x[26] & ~x[30] & ~x[42] & ~x[43] & ~x[58] & ~x[61];
			partial_clause[241] 	= 1'b1;
			partial_clause[242] 	= ~x[6] & ~x[9] & ~x[18] & ~x[24] & ~x[29] & ~x[30] & ~x[40] & ~x[50] & ~x[59] & ~x[61] & ~x[63];
			partial_clause[243] 	= ~x[0] & ~x[1] & ~x[2] & ~x[13] & ~x[15] & ~x[29] & ~x[32] & ~x[39] & ~x[43] & ~x[50] & ~x[57];
			partial_clause[244] 	= ~x[40];
			partial_clause[245] 	= 1'b1;
			partial_clause[246] 	= ~x[27];
			partial_clause[247] 	= ~x[2] & ~x[5] & ~x[6] & ~x[10] & ~x[15] & ~x[17] & ~x[19] & ~x[20] & ~x[23] & ~x[26] & ~x[32] & ~x[34] & ~x[38] & ~x[40] & ~x[42] & ~x[49] & ~x[50] & ~x[52] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[248] 	= ~x[1] & ~x[5] & ~x[10] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[21] & ~x[23] & ~x[24] & ~x[28] & ~x[31] & ~x[46] & ~x[48] & ~x[51] & ~x[52];
			partial_clause[249] 	= ~x[24] & ~x[43] & ~x[48];
			partial_clause[250] 	= ~x[4] & ~x[9] & ~x[10] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[24] & ~x[25] & ~x[27] & ~x[28] & ~x[36] & ~x[38] & ~x[39] & ~x[41] & ~x[42] & ~x[43] & ~x[47] & ~x[48] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[59] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[251] 	= ~x[3];
			partial_clause[252] 	= ~x[5] & ~x[11] & ~x[19] & ~x[22] & ~x[23] & ~x[26] & ~x[33] & ~x[34] & ~x[35] & ~x[41] & ~x[42] & ~x[44] & ~x[45] & ~x[46] & ~x[49] & ~x[52] & ~x[53] & ~x[54] & ~x[57] & ~x[58] & ~x[61];
			partial_clause[253] 	= 1'b1;
			partial_clause[254] 	= ~x[10] & ~x[19] & ~x[24] & ~x[25] & ~x[34] & ~x[40];
			partial_clause[255] 	= ~x[5] & ~x[22] & ~x[30] & ~x[63];
			partial_clause[256] 	= 1'b1;
			partial_clause[257] 	= ~x[38] & ~x[46];
			partial_clause[258] 	= ~x[5] & ~x[10] & ~x[25] & ~x[61];
			partial_clause[259] 	= 1'b1;
			partial_clause[260] 	= ~x[2] & ~x[33] & ~x[44] & ~x[61];
			partial_clause[261] 	= ~x[18] & ~x[19] & ~x[23] & ~x[29] & ~x[30] & ~x[36] & ~x[42] & ~x[45] & ~x[48] & ~x[49] & ~x[59];
			partial_clause[262] 	= ~x[31] & ~x[33];
			partial_clause[263] 	= ~x[53];
			partial_clause[264] 	= ~x[56] & ~x[59];
			partial_clause[265] 	= 1'b1;
			partial_clause[266] 	= ~x[0] & ~x[1] & ~x[5] & ~x[7] & ~x[10] & ~x[13] & ~x[24] & ~x[31] & ~x[32] & ~x[40] & ~x[43] & ~x[53] & ~x[56];
			partial_clause[267] 	= ~x[0] & ~x[1] & ~x[2] & ~x[5] & ~x[10] & ~x[17] & ~x[18] & ~x[23] & ~x[28] & ~x[29] & ~x[30] & ~x[33] & ~x[38] & ~x[52] & ~x[57] & ~x[60] & ~x[61];
			partial_clause[268] 	= ~x[6] & ~x[8] & ~x[22] & ~x[29] & ~x[32] & ~x[36] & ~x[38] & ~x[40] & ~x[44] & ~x[46] & ~x[49] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[62];
			partial_clause[269] 	= ~x[2] & ~x[6] & ~x[8] & ~x[13] & ~x[14] & ~x[15] & ~x[17] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[24] & ~x[25] & ~x[26] & ~x[29] & ~x[30] & ~x[32] & ~x[36] & ~x[38] & ~x[39] & ~x[40] & ~x[41] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[54] & ~x[56] & ~x[59] & ~x[60];
			partial_clause[270] 	= 1'b1;
			partial_clause[271] 	= ~x[15] & ~x[20];
			partial_clause[272] 	= ~x[1] & ~x[11] & ~x[12] & ~x[13] & ~x[21] & ~x[25] & ~x[29] & ~x[30] & ~x[31] & ~x[41] & ~x[49] & ~x[55] & ~x[60];
			partial_clause[273] 	= ~x[2] & ~x[7] & ~x[8] & ~x[14] & ~x[15] & ~x[21] & ~x[23] & ~x[27] & ~x[29] & ~x[31] & ~x[32] & ~x[33] & ~x[34] & ~x[35] & ~x[39] & ~x[40] & ~x[42] & ~x[43] & ~x[44] & ~x[49] & ~x[51] & ~x[55] & ~x[56] & ~x[63];
			partial_clause[274] 	= ~x[9] & ~x[14] & ~x[20] & ~x[25] & ~x[27] & ~x[34] & ~x[41] & ~x[48] & ~x[54];
			partial_clause[275] 	= ~x[12] & ~x[22] & ~x[40] & ~x[54];
			partial_clause[276] 	= ~x[21] & ~x[22] & ~x[26] & ~x[33] & ~x[35] & ~x[39] & ~x[63];
			partial_clause[277] 	= ~x[2] & ~x[30] & ~x[41] & ~x[47] & ~x[61] & ~x[62];
			partial_clause[278] 	= 1'b1;
			partial_clause[279] 	= ~x[4] & ~x[5] & ~x[6] & ~x[13] & ~x[14] & ~x[16] & ~x[17] & ~x[22] & ~x[23] & ~x[30] & ~x[45] & ~x[52] & ~x[53] & ~x[54] & ~x[56] & ~x[57] & ~x[58] & ~x[59] & ~x[60];
			partial_clause[280] 	= 1'b1;
			partial_clause[281] 	= ~x[4] & ~x[5] & ~x[28] & ~x[40] & ~x[43] & ~x[53] & ~x[57] & ~x[63];
			partial_clause[282] 	= ~x[26] & ~x[29] & ~x[50];
			partial_clause[283] 	= ~x[28] & ~x[58];
			partial_clause[284] 	= ~x[16] & ~x[18] & ~x[32] & ~x[63];
			partial_clause[285] 	= ~x[4];
			partial_clause[286] 	= ~x[19] & ~x[36] & ~x[37];
			partial_clause[287] 	= ~x[0] & ~x[3] & ~x[7] & ~x[9] & ~x[19] & ~x[20] & ~x[23] & ~x[25] & ~x[26] & ~x[31] & ~x[32] & ~x[41] & ~x[44] & ~x[51] & ~x[55] & ~x[56] & ~x[59];
			partial_clause[288] 	= ~x[18] & ~x[21];
			partial_clause[289] 	= ~x[4] & ~x[6] & ~x[19] & ~x[20] & ~x[54] & ~x[60] & ~x[63];
			partial_clause[290] 	= ~x[22] & ~x[46] & ~x[51];
			partial_clause[291] 	= ~x[52] & ~x[57];
			partial_clause[292] 	= ~x[28];
			partial_clause[293] 	= ~x[2] & ~x[50] & ~x[51] & ~x[55];
			partial_clause[294] 	= ~x[12] & ~x[26] & ~x[40];
			partial_clause[295] 	= ~x[58];
			partial_clause[296] 	= 1'b1;
			partial_clause[297] 	= ~x[15] & ~x[34] & ~x[42] & ~x[54] & ~x[62] & ~x[63];
			partial_clause[298] 	= 1'b1;
			partial_clause[299] 	= ~x[19] & ~x[22] & ~x[34] & ~x[40] & ~x[52] & ~x[55] & ~x[62];
			partial_clause[300] 	= ~x[25] & ~x[46] & ~x[54] & ~x[56] & ~x[58];
			partial_clause[301] 	= ~x[9] & ~x[18] & ~x[46] & ~x[48] & ~x[50];
			partial_clause[302] 	= ~x[3] & ~x[32];
			partial_clause[303] 	= ~x[3] & ~x[16] & ~x[33] & ~x[47];
			partial_clause[304] 	= ~x[25];
			partial_clause[305] 	= ~x[0] & ~x[13] & ~x[37] & ~x[62];
			partial_clause[306] 	= ~x[10] & ~x[14] & ~x[23] & ~x[26] & ~x[35] & ~x[41] & ~x[48] & ~x[54];
			partial_clause[307] 	= ~x[21] & ~x[35] & ~x[46] & ~x[47] & ~x[49] & ~x[53] & ~x[54] & ~x[57] & ~x[62];
			partial_clause[308] 	= ~x[7] & ~x[11] & ~x[15] & ~x[21] & ~x[23] & ~x[29] & ~x[30] & ~x[35] & ~x[40] & ~x[51] & ~x[56] & ~x[60];
			partial_clause[309] 	= ~x[3] & ~x[12] & ~x[14] & ~x[46] & ~x[47] & ~x[55];
			partial_clause[310] 	= 1'b1;
			partial_clause[311] 	= ~x[19] & ~x[20] & ~x[32] & ~x[35] & ~x[37] & ~x[41] & ~x[48] & ~x[50] & ~x[55] & ~x[59];
			partial_clause[312] 	= 1'b1;
			partial_clause[313] 	= ~x[52] & ~x[59];
			partial_clause[314] 	= ~x[9] & ~x[19];
			partial_clause[315] 	= ~x[14] & ~x[53] & ~x[63];
			partial_clause[316] 	= ~x[6] & ~x[7] & ~x[9] & ~x[14] & ~x[18] & ~x[27] & ~x[29] & ~x[39] & ~x[42] & ~x[44] & ~x[50] & ~x[62];
			partial_clause[317] 	= ~x[15] & ~x[16] & ~x[36] & ~x[38] & ~x[47] & ~x[60];
			partial_clause[318] 	= ~x[0] & ~x[11] & ~x[33] & ~x[47];
			partial_clause[319] 	= ~x[56];
			partial_clause[320] 	= ~x[10] & ~x[13] & ~x[17] & ~x[23] & ~x[45] & ~x[49] & ~x[52] & ~x[55];
			partial_clause[321] 	= ~x[0] & ~x[1] & ~x[8] & ~x[10] & ~x[15] & ~x[18] & ~x[27] & ~x[34] & ~x[48] & ~x[49] & ~x[53];
			partial_clause[322] 	= ~x[47] & ~x[61] & ~x[62];
			partial_clause[323] 	= ~x[11] & ~x[60];
			partial_clause[324] 	= ~x[8] & ~x[11] & ~x[17] & ~x[59] & ~x[60];
			partial_clause[325] 	= ~x[3] & ~x[8] & ~x[10] & ~x[11] & ~x[14] & ~x[16] & ~x[17] & ~x[19] & ~x[20] & ~x[23] & ~x[24] & ~x[26] & ~x[27] & ~x[30] & ~x[31] & ~x[33] & ~x[34] & ~x[36] & ~x[37] & ~x[38] & ~x[41] & ~x[42] & ~x[43] & ~x[49] & ~x[51] & ~x[54] & ~x[58] & ~x[59] & ~x[62] & ~x[63];
			partial_clause[326] 	= ~x[0] & ~x[3] & ~x[8] & ~x[11] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[19] & ~x[20] & ~x[28] & ~x[41] & ~x[47] & ~x[49] & ~x[51] & ~x[52] & ~x[61] & ~x[63];
			partial_clause[327] 	= ~x[16] & ~x[21] & ~x[26] & ~x[50] & ~x[58];
			partial_clause[328] 	= ~x[20] & ~x[47] & ~x[57] & ~x[60] & ~x[61];
			partial_clause[329] 	= 1'b1;
			partial_clause[330] 	= ~x[19] & ~x[26] & ~x[29] & ~x[36];
			partial_clause[331] 	= ~x[1] & ~x[61];
			partial_clause[332] 	= ~x[39] & ~x[56] & ~x[61];
			partial_clause[333] 	= ~x[14] & ~x[43];
			partial_clause[334] 	= ~x[1] & ~x[9];
			partial_clause[335] 	= ~x[24] & ~x[29] & ~x[30];
			partial_clause[336] 	= 1'b1;
			partial_clause[337] 	= ~x[0] & ~x[3] & ~x[7] & ~x[12] & ~x[16] & ~x[19] & ~x[23] & ~x[38] & ~x[43] & ~x[46] & ~x[47] & ~x[49] & ~x[62];
			partial_clause[338] 	= 1'b1;
			partial_clause[339] 	= ~x[0] & ~x[4] & ~x[11] & ~x[14] & ~x[15] & ~x[27] & ~x[29] & ~x[33] & ~x[34] & ~x[38] & ~x[39] & ~x[42] & ~x[47] & ~x[55] & ~x[57] & ~x[60];
			partial_clause[340] 	= ~x[6] & ~x[9] & ~x[11] & ~x[13] & ~x[14] & ~x[16] & ~x[32] & ~x[33] & ~x[41] & ~x[44] & ~x[47] & ~x[50] & ~x[54] & ~x[58];
			partial_clause[341] 	= 1'b1;
			partial_clause[342] 	= ~x[4] & ~x[19] & ~x[25] & ~x[31] & ~x[32] & ~x[36] & ~x[40] & ~x[41] & ~x[42] & ~x[45] & ~x[51] & ~x[54] & ~x[55] & ~x[56] & ~x[61];
			partial_clause[343] 	= ~x[14] & ~x[15] & ~x[27] & ~x[30] & ~x[32] & ~x[52] & ~x[53] & ~x[61] & ~x[63];
			partial_clause[344] 	= ~x[1] & ~x[7] & ~x[22] & ~x[23] & ~x[25] & ~x[36] & ~x[44] & ~x[50] & ~x[51];
			partial_clause[345] 	= ~x[37] & ~x[43] & ~x[56];
			partial_clause[346] 	= ~x[3] & ~x[13] & ~x[16] & ~x[17];
			partial_clause[347] 	= ~x[0] & ~x[1] & ~x[13] & ~x[15] & ~x[40] & ~x[45] & ~x[55];
			partial_clause[348] 	= ~x[12] & ~x[40];
			partial_clause[349] 	= ~x[48] & ~x[62];
			partial_clause[350] 	= ~x[0] & ~x[1] & ~x[2] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[12] & ~x[15] & ~x[19] & ~x[21] & ~x[23] & ~x[24] & ~x[26] & ~x[28] & ~x[29] & ~x[33] & ~x[34] & ~x[36] & ~x[37] & ~x[42] & ~x[44] & ~x[45] & ~x[48] & ~x[51] & ~x[53] & ~x[56] & ~x[58] & ~x[61];
			partial_clause[351] 	= 1'b1;
			partial_clause[352] 	= 1'b1;
			partial_clause[353] 	= ~x[0] & ~x[5] & ~x[13] & ~x[20] & ~x[52] & ~x[61];
			partial_clause[354] 	= ~x[14] & ~x[21] & ~x[26] & ~x[28] & ~x[30] & ~x[41] & ~x[42];
			partial_clause[355] 	= ~x[2] & ~x[12] & ~x[22] & ~x[50] & ~x[55];
			partial_clause[356] 	= ~x[9] & ~x[10] & ~x[21] & ~x[61];
			partial_clause[357] 	= 1'b1;
			partial_clause[358] 	= ~x[2] & ~x[13] & ~x[23] & ~x[26] & ~x[31] & ~x[42] & ~x[49] & ~x[52] & ~x[53] & ~x[60] & ~x[62];
			partial_clause[359] 	= ~x[2] & ~x[3] & ~x[7] & ~x[13] & ~x[16] & ~x[17] & ~x[33] & ~x[39] & ~x[40];
			partial_clause[360] 	= ~x[0] & ~x[3] & ~x[4] & ~x[5] & ~x[9] & ~x[10] & ~x[11] & ~x[17] & ~x[21] & ~x[24] & ~x[26] & ~x[28] & ~x[30] & ~x[33] & ~x[38] & ~x[44] & ~x[46] & ~x[50] & ~x[51] & ~x[53] & ~x[56] & ~x[57] & ~x[58] & ~x[62];
			partial_clause[361] 	= ~x[10] & ~x[11] & ~x[21] & ~x[24] & ~x[30] & ~x[32] & ~x[35] & ~x[39] & ~x[44] & ~x[46] & ~x[52] & ~x[53] & ~x[54];
			partial_clause[362] 	= ~x[14] & ~x[23] & ~x[29] & ~x[34] & ~x[37] & ~x[38] & ~x[49] & ~x[53] & ~x[56] & ~x[58];
			partial_clause[363] 	= ~x[2] & ~x[9] & ~x[16] & ~x[23] & ~x[25] & ~x[27] & ~x[30] & ~x[38] & ~x[40] & ~x[43] & ~x[53] & ~x[57];
			partial_clause[364] 	= ~x[1] & ~x[11] & ~x[12] & ~x[30] & ~x[49] & ~x[51] & ~x[55] & ~x[59];
			partial_clause[365] 	= ~x[8] & ~x[11] & ~x[59];
			partial_clause[366] 	= ~x[3] & ~x[4] & ~x[8] & ~x[10] & ~x[15] & ~x[32] & ~x[34] & ~x[36] & ~x[39] & ~x[50] & ~x[52] & ~x[54] & ~x[57] & ~x[61];
			partial_clause[367] 	= ~x[0] & ~x[10] & ~x[17] & ~x[18] & ~x[26] & ~x[37] & ~x[46] & ~x[56] & ~x[57] & ~x[62];
			partial_clause[368] 	= 1'b1;
			partial_clause[369] 	= ~x[18] & ~x[50] & ~x[51];
			partial_clause[370] 	= ~x[4] & ~x[17] & ~x[20] & ~x[24] & ~x[29] & ~x[34] & ~x[60];
			partial_clause[371] 	= ~x[1];
			partial_clause[372] 	= ~x[18] & ~x[26] & ~x[27] & ~x[58] & ~x[60];
			partial_clause[373] 	= 1'b1;
			partial_clause[374] 	= ~x[4] & ~x[36] & ~x[45] & ~x[54];
			partial_clause[375] 	= ~x[18];
			partial_clause[376] 	= ~x[4] & ~x[12] & ~x[15] & ~x[24] & ~x[28] & ~x[30] & ~x[32] & ~x[40] & ~x[42] & ~x[44] & ~x[46] & ~x[55];
			partial_clause[377] 	= ~x[9] & ~x[19] & ~x[22] & ~x[23] & ~x[25] & ~x[40] & ~x[42] & ~x[52] & ~x[59];
			partial_clause[378] 	= ~x[1];
			partial_clause[379] 	= ~x[1] & ~x[20] & ~x[24] & ~x[35] & ~x[43] & ~x[46] & ~x[56] & ~x[62];
			partial_clause[380] 	= 1'b1;
			partial_clause[381] 	= ~x[1] & ~x[3] & ~x[4] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[26] & ~x[27] & ~x[29] & ~x[37] & ~x[44] & ~x[50] & ~x[52] & ~x[54] & ~x[56];
			partial_clause[382] 	= 1'b1;
			partial_clause[383] 	= 1'b1;
			partial_clause[384] 	= 1'b1;
			partial_clause[385] 	= 1'b1;
			partial_clause[386] 	= ~x[37] & ~x[52] & ~x[57];
			partial_clause[387] 	= ~x[3] & ~x[6] & ~x[8] & ~x[12] & ~x[13] & ~x[19] & ~x[28] & ~x[33] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[44] & ~x[48] & ~x[50] & ~x[60] & ~x[62];
			partial_clause[388] 	= ~x[2] & ~x[3] & ~x[7] & ~x[9] & ~x[13] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[20] & ~x[21] & ~x[22] & ~x[25] & ~x[29] & ~x[36] & ~x[38] & ~x[46] & ~x[49] & ~x[51] & ~x[53] & ~x[54] & ~x[59] & ~x[63];
			partial_clause[389] 	= 1'b1;
			partial_clause[390] 	= ~x[2] & ~x[6] & ~x[9] & ~x[13] & ~x[15] & ~x[17] & ~x[30] & ~x[31] & ~x[32] & ~x[39] & ~x[45] & ~x[50] & ~x[57];
			partial_clause[391] 	= 1'b1;
			partial_clause[392] 	= 1'b1;
			partial_clause[393] 	= 1'b1;
			partial_clause[394] 	= ~x[9] & ~x[28] & ~x[49] & ~x[50] & ~x[53] & ~x[56];
			partial_clause[395] 	= 1'b1;
			partial_clause[396] 	= 1'b1;
			partial_clause[397] 	= 1'b1;
			partial_clause[398] 	= ~x[14];
			partial_clause[399] 	= 1'b1;
			partial_clause[400] 	= ~x[0] & ~x[6] & ~x[8] & ~x[14] & ~x[15] & ~x[19] & ~x[26] & ~x[41] & ~x[52] & ~x[53];
			partial_clause[401] 	= ~x[3] & ~x[6] & ~x[10] & ~x[13] & ~x[16] & ~x[18] & ~x[22] & ~x[23] & ~x[24] & ~x[29] & ~x[33] & ~x[34] & ~x[42] & ~x[43] & ~x[45] & ~x[47] & ~x[56] & ~x[57] & ~x[58];
			partial_clause[402] 	= ~x[3] & ~x[4] & ~x[6] & ~x[10] & ~x[23] & ~x[25] & ~x[34] & ~x[44] & ~x[53] & ~x[55] & ~x[60];
			partial_clause[403] 	= ~x[3] & ~x[56];
			partial_clause[404] 	= 1'b1;
			partial_clause[405] 	= ~x[5] & ~x[10] & ~x[21] & ~x[22] & ~x[44] & ~x[53] & ~x[59];
			partial_clause[406] 	= ~x[13] & ~x[15] & ~x[38] & ~x[54] & ~x[56];
			partial_clause[407] 	= ~x[8];
			partial_clause[408] 	= ~x[3] & ~x[21] & ~x[31] & ~x[38] & ~x[43] & ~x[46] & ~x[51];
			partial_clause[409] 	= ~x[6] & ~x[13] & ~x[14] & ~x[18] & ~x[21] & ~x[25] & ~x[27] & ~x[28] & ~x[30] & ~x[43] & ~x[44] & ~x[46] & ~x[49] & ~x[51] & ~x[52] & ~x[56] & ~x[58] & ~x[60] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[410] 	= ~x[2] & ~x[12] & ~x[33] & ~x[35] & ~x[42] & ~x[43] & ~x[51] & ~x[61];
			partial_clause[411] 	= ~x[11] & ~x[23] & ~x[40] & ~x[45] & ~x[56] & ~x[61];
			partial_clause[412] 	= ~x[0] & ~x[1] & ~x[4] & ~x[5] & ~x[8] & ~x[9] & ~x[24] & ~x[29] & ~x[32] & ~x[36] & ~x[41] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[53] & ~x[54] & ~x[55] & ~x[58] & ~x[62];
			partial_clause[413] 	= ~x[9] & ~x[11] & ~x[18] & ~x[29] & ~x[38] & ~x[52];
			partial_clause[414] 	= ~x[3] & ~x[24] & ~x[27] & ~x[32] & ~x[38] & ~x[47] & ~x[48];
			partial_clause[415] 	= ~x[1] & ~x[5] & ~x[7] & ~x[10] & ~x[12] & ~x[28] & ~x[34] & ~x[45] & ~x[46];
			partial_clause[416] 	= ~x[2] & ~x[8] & ~x[9] & ~x[15] & ~x[21] & ~x[31] & ~x[36] & ~x[39] & ~x[44] & ~x[45] & ~x[48] & ~x[49] & ~x[53] & ~x[54] & ~x[60] & ~x[61];
			partial_clause[417] 	= ~x[2] & ~x[21] & ~x[22] & ~x[39];
			partial_clause[418] 	= ~x[4] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[23] & ~x[25] & ~x[33] & ~x[34] & ~x[35] & ~x[36] & ~x[40] & ~x[41] & ~x[49] & ~x[57] & ~x[60] & ~x[61];
			partial_clause[419] 	= 1'b1;
			partial_clause[420] 	= 1'b1;
			partial_clause[421] 	= ~x[26] & ~x[36] & ~x[40] & ~x[47] & ~x[48] & ~x[57] & ~x[60];
			partial_clause[422] 	= ~x[19] & ~x[29] & ~x[43] & ~x[47] & ~x[48] & ~x[58] & ~x[62];
			partial_clause[423] 	= ~x[9] & ~x[17] & ~x[25] & ~x[29] & ~x[45] & ~x[63];
			partial_clause[424] 	= ~x[15] & ~x[19] & ~x[30] & ~x[31] & ~x[41] & ~x[46] & ~x[52];
			partial_clause[425] 	= ~x[32] & ~x[35];
			partial_clause[426] 	= ~x[0] & ~x[6] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[20] & ~x[21] & ~x[24] & ~x[26] & ~x[27] & ~x[28] & ~x[30] & ~x[38] & ~x[41] & ~x[51] & ~x[52] & ~x[55] & ~x[59] & ~x[63];
			partial_clause[427] 	= ~x[9] & ~x[23] & ~x[28] & ~x[29] & ~x[36] & ~x[38] & ~x[39] & ~x[44] & ~x[47] & ~x[59];
			partial_clause[428] 	= ~x[11];
			partial_clause[429] 	= 1'b1;
			partial_clause[430] 	= ~x[3] & ~x[4] & ~x[5] & ~x[8] & ~x[12] & ~x[18] & ~x[20] & ~x[24] & ~x[25] & ~x[26] & ~x[29] & ~x[33] & ~x[35] & ~x[37] & ~x[38] & ~x[43] & ~x[46] & ~x[48] & ~x[51] & ~x[54] & ~x[55];
			partial_clause[431] 	= ~x[7] & ~x[15] & ~x[39] & ~x[44];
			partial_clause[432] 	= ~x[4] & ~x[5] & ~x[14] & ~x[15] & ~x[21] & ~x[30] & ~x[36] & ~x[40] & ~x[48] & ~x[55] & ~x[57] & ~x[62];
			partial_clause[433] 	= ~x[21] & ~x[29] & ~x[46];
			partial_clause[434] 	= ~x[12] & ~x[26] & ~x[53];
			partial_clause[435] 	= ~x[1] & ~x[6] & ~x[7] & ~x[16] & ~x[17] & ~x[24] & ~x[25] & ~x[30] & ~x[34] & ~x[35] & ~x[39] & ~x[40] & ~x[41] & ~x[48] & ~x[49] & ~x[54] & ~x[55] & ~x[63];
			partial_clause[436] 	= ~x[0] & ~x[1] & ~x[11] & ~x[22] & ~x[25] & ~x[31] & ~x[33] & ~x[37] & ~x[40] & ~x[47] & ~x[50] & ~x[54] & ~x[60];
			partial_clause[437] 	= ~x[1] & ~x[3] & ~x[4] & ~x[8] & ~x[13] & ~x[15] & ~x[25] & ~x[26] & ~x[27] & ~x[36] & ~x[37] & ~x[39] & ~x[45] & ~x[48] & ~x[52] & ~x[55] & ~x[58];
			partial_clause[438] 	= 1'b1;
			partial_clause[439] 	= ~x[4] & ~x[5] & ~x[15] & ~x[16] & ~x[21] & ~x[57];
			partial_clause[440] 	= ~x[29] & ~x[36];
			partial_clause[441] 	= ~x[8] & ~x[10] & ~x[12] & ~x[18] & ~x[19];
			partial_clause[442] 	= 1'b1;
			partial_clause[443] 	= ~x[2] & ~x[5] & ~x[9] & ~x[13] & ~x[14] & ~x[19] & ~x[20] & ~x[22] & ~x[28] & ~x[36] & ~x[43] & ~x[48] & ~x[52] & ~x[55] & ~x[62];
			partial_clause[444] 	= 1'b1;
			partial_clause[445] 	= ~x[45];
			partial_clause[446] 	= ~x[0] & ~x[2] & ~x[4] & ~x[5] & ~x[15] & ~x[18] & ~x[34] & ~x[47] & ~x[55] & ~x[57];
			partial_clause[447] 	= ~x[0] & ~x[1] & ~x[5] & ~x[10] & ~x[14] & ~x[20] & ~x[24] & ~x[25] & ~x[30];
			partial_clause[448] 	= 1'b1;
			partial_clause[449] 	= ~x[6] & ~x[16] & ~x[22] & ~x[25] & ~x[32] & ~x[35] & ~x[36] & ~x[39] & ~x[41] & ~x[42] & ~x[51] & ~x[59];
			partial_clause[450] 	= ~x[6] & ~x[8] & ~x[33] & ~x[47] & ~x[51] & ~x[56];
			partial_clause[451] 	= 1'b1;
			partial_clause[452] 	= ~x[26] & ~x[45];
			partial_clause[453] 	= ~x[10] & ~x[61];
			partial_clause[454] 	= ~x[3] & ~x[8] & ~x[49];
			partial_clause[455] 	= ~x[2] & ~x[17] & ~x[20] & ~x[28] & ~x[63];
			partial_clause[456] 	= ~x[0] & ~x[10] & ~x[19] & ~x[21] & ~x[26] & ~x[33] & ~x[37] & ~x[43] & ~x[46] & ~x[47] & ~x[48];
			partial_clause[457] 	= ~x[12] & ~x[20];
			partial_clause[458] 	= ~x[4] & ~x[8] & ~x[12] & ~x[23] & ~x[33] & ~x[34] & ~x[41] & ~x[42] & ~x[44] & ~x[46] & ~x[47] & ~x[54];
			partial_clause[459] 	= ~x[2] & ~x[16] & ~x[18] & ~x[26] & ~x[29] & ~x[33] & ~x[43] & ~x[48] & ~x[54] & ~x[59];
			partial_clause[460] 	= ~x[4] & ~x[6] & ~x[13] & ~x[15] & ~x[29] & ~x[30] & ~x[32] & ~x[37] & ~x[43] & ~x[45] & ~x[47] & ~x[50] & ~x[56] & ~x[57];
			partial_clause[461] 	= ~x[19] & ~x[20] & ~x[24] & ~x[28] & ~x[32] & ~x[35] & ~x[36] & ~x[37] & ~x[50] & ~x[51] & ~x[57] & ~x[59];
			partial_clause[462] 	= ~x[51];
			partial_clause[463] 	= 1'b1;
			partial_clause[464] 	= ~x[16] & ~x[18];
			partial_clause[465] 	= ~x[20] & ~x[26] & ~x[30] & ~x[31] & ~x[32] & ~x[34] & ~x[38] & ~x[41] & ~x[55] & ~x[58] & ~x[61];
			partial_clause[466] 	= ~x[3] & ~x[4] & ~x[7] & ~x[10] & ~x[11] & ~x[13] & ~x[16] & ~x[18] & ~x[24] & ~x[32] & ~x[36] & ~x[39] & ~x[41] & ~x[43] & ~x[53] & ~x[57] & ~x[59] & ~x[62];
			partial_clause[467] 	= ~x[7] & ~x[46] & ~x[52] & ~x[61];
			partial_clause[468] 	= ~x[7] & ~x[15] & ~x[18] & ~x[29] & ~x[54] & ~x[57];
			partial_clause[469] 	= ~x[2] & ~x[4] & ~x[10] & ~x[11] & ~x[22] & ~x[29] & ~x[32] & ~x[38] & ~x[39] & ~x[40] & ~x[46];
			partial_clause[470] 	= ~x[49];
			partial_clause[471] 	= ~x[18] & ~x[22] & ~x[31] & ~x[37] & ~x[38] & ~x[42] & ~x[48] & ~x[51] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[59] & ~x[60];
			partial_clause[472] 	= ~x[3] & ~x[35] & ~x[47];
			partial_clause[473] 	= ~x[1] & ~x[2] & ~x[3] & ~x[9] & ~x[12] & ~x[16] & ~x[17] & ~x[42] & ~x[45] & ~x[46];
			partial_clause[474] 	= 1'b1;
			partial_clause[475] 	= ~x[3] & ~x[11] & ~x[14] & ~x[18] & ~x[22] & ~x[24] & ~x[27] & ~x[41] & ~x[57];
			partial_clause[476] 	= ~x[50];
			partial_clause[477] 	= ~x[2] & ~x[3] & ~x[7] & ~x[10] & ~x[15] & ~x[20] & ~x[23] & ~x[24] & ~x[42] & ~x[50] & ~x[57] & ~x[59] & ~x[63];
			partial_clause[478] 	= ~x[0] & ~x[7] & ~x[11] & ~x[18] & ~x[19] & ~x[35] & ~x[36] & ~x[38] & ~x[39] & ~x[43] & ~x[45] & ~x[46] & ~x[52] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[63];
			partial_clause[479] 	= 1'b1;
			partial_clause[480] 	= ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[8] & ~x[10] & ~x[11] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[25] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & ~x[31] & ~x[32] & ~x[33] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[38] & ~x[39] & ~x[41] & ~x[45] & ~x[46] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[59] & ~x[60] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[481] 	= ~x[19] & ~x[36] & ~x[53] & ~x[57];
			partial_clause[482] 	= ~x[19];
			partial_clause[483] 	= ~x[3] & ~x[38] & ~x[40] & ~x[52];
			partial_clause[484] 	= ~x[23] & ~x[38] & ~x[44];
			partial_clause[485] 	= 1'b1;
			partial_clause[486] 	= ~x[0] & ~x[1] & ~x[12] & ~x[23] & ~x[30] & ~x[43] & ~x[57] & ~x[61];
			partial_clause[487] 	= ~x[4] & ~x[7] & ~x[13] & ~x[17] & ~x[33] & ~x[36] & ~x[40] & ~x[51] & ~x[62];
			partial_clause[488] 	= 1'b1;
			partial_clause[489] 	= 1'b1;
			partial_clause[490] 	= 1'b1;
			partial_clause[491] 	= ~x[32] & ~x[41] & ~x[43] & ~x[46] & ~x[50];
			partial_clause[492] 	= ~x[2] & ~x[6] & ~x[9] & ~x[15] & ~x[25] & ~x[43] & ~x[53] & ~x[55] & ~x[61];
			partial_clause[493] 	= ~x[8];
			partial_clause[494] 	= ~x[7] & ~x[25] & ~x[28] & ~x[50];
			partial_clause[495] 	= ~x[2] & ~x[3] & ~x[5] & ~x[7] & ~x[14] & ~x[28] & ~x[29] & ~x[43] & ~x[45] & ~x[49] & ~x[50] & ~x[58];
			partial_clause[496] 	= 1'b1;
			partial_clause[497] 	= ~x[60];
			partial_clause[498] 	= 1'b1;
			partial_clause[499] 	= ~x[5] & ~x[17] & ~x[27] & ~x[37] & ~x[43] & ~x[52];
		end
	end
endmodule


module HCB_1 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[0] & ~x[1] & ~x[3] & ~x[5] & ~x[7] & ~x[9] & ~x[10] & ~x[13] & ~x[14] & ~x[16] & ~x[23] & ~x[28] & ~x[32] & ~x[33] & ~x[39] & ~x[40] & ~x[42] & ~x[44] & ~x[46] & ~x[48] & ~x[49] & ~x[52] & ~x[57];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[4] & ~x[9] & ~x[11] & ~x[12] & ~x[19] & ~x[42] & ~x[63];
			partial_clause[2] 	= partial_clause_prev[2] & 1'b1;
			partial_clause[3] 	= partial_clause_prev[3] & ~x[12] & ~x[18] & ~x[34] & ~x[35] & ~x[52];
			partial_clause[4] 	= partial_clause_prev[4] & ~x[33] & ~x[45] & ~x[55];
			partial_clause[5] 	= partial_clause_prev[5] & ~x[4] & ~x[5] & ~x[6] & ~x[15] & ~x[21] & ~x[22] & ~x[24] & ~x[27] & ~x[29] & ~x[30] & ~x[33] & ~x[37] & ~x[38] & ~x[46] & ~x[58];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[14] & ~x[26] & ~x[43] & ~x[46];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[2] & ~x[4] & ~x[8] & ~x[26] & ~x[27] & ~x[28] & ~x[41] & ~x[45] & ~x[46] & ~x[55] & ~x[56];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[1] & ~x[3] & ~x[6] & ~x[9] & ~x[12] & ~x[18] & ~x[23] & ~x[24] & ~x[25] & ~x[27] & ~x[38] & ~x[43] & ~x[46] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[56] & ~x[58];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[5] & ~x[6] & ~x[9] & ~x[11] & ~x[14] & ~x[17] & ~x[18] & ~x[30] & ~x[32] & ~x[33] & ~x[47] & ~x[53] & ~x[56] & ~x[57] & ~x[58] & ~x[59];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[15] & ~x[20] & ~x[24] & ~x[27] & ~x[35] & ~x[49] & ~x[53] & ~x[54] & ~x[57];
			partial_clause[11] 	= partial_clause_prev[11] & ~x[2] & ~x[14] & ~x[21] & ~x[22] & ~x[33] & ~x[41] & ~x[47] & ~x[49] & ~x[56] & ~x[57];
			partial_clause[12] 	= partial_clause_prev[12] & ~x[14] & ~x[16] & ~x[17] & ~x[21] & ~x[22] & ~x[24] & ~x[26] & ~x[28] & ~x[30] & ~x[40] & ~x[47] & ~x[51] & ~x[53] & ~x[56] & ~x[60];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[2] & ~x[3] & ~x[7] & ~x[8] & ~x[10] & ~x[17] & ~x[23] & ~x[27] & ~x[30] & ~x[43] & ~x[46] & ~x[48] & ~x[49] & ~x[57];
			partial_clause[14] 	= partial_clause_prev[14] & 1'b1;
			partial_clause[15] 	= partial_clause_prev[15] & 1'b1;
			partial_clause[16] 	= partial_clause_prev[16] & ~x[0] & ~x[33] & ~x[41] & ~x[42] & ~x[49] & ~x[52] & ~x[54];
			partial_clause[17] 	= partial_clause_prev[17] & 1'b1;
			partial_clause[18] 	= partial_clause_prev[18] & ~x[4] & ~x[21] & ~x[24];
			partial_clause[19] 	= partial_clause_prev[19] & ~x[9] & ~x[13] & ~x[17] & ~x[18] & ~x[22] & ~x[47] & ~x[48];
			partial_clause[20] 	= partial_clause_prev[20] & ~x[15] & ~x[29] & ~x[38] & ~x[44];
			partial_clause[21] 	= partial_clause_prev[21] & ~x[5] & ~x[25];
			partial_clause[22] 	= partial_clause_prev[22] & ~x[1] & ~x[23] & ~x[28] & ~x[30];
			partial_clause[23] 	= partial_clause_prev[23] & ~x[7] & ~x[10] & ~x[12] & ~x[14] & ~x[15] & ~x[16] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[25] & ~x[26] & ~x[38] & ~x[39] & ~x[40] & ~x[41] & ~x[43] & ~x[45] & ~x[46] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[0] & ~x[1] & ~x[2] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[15] & ~x[16] & ~x[17] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[27] & ~x[29] & ~x[36] & ~x[40] & ~x[44] & ~x[47] & ~x[50] & ~x[51] & ~x[52] & ~x[54] & ~x[55] & ~x[56];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[0] & ~x[2] & ~x[6] & ~x[9] & ~x[10] & ~x[13] & ~x[14] & ~x[17] & ~x[18] & ~x[20] & ~x[23] & ~x[25] & ~x[27] & ~x[28] & ~x[30] & ~x[31] & ~x[32] & ~x[39] & ~x[41] & ~x[42] & ~x[43] & ~x[45] & ~x[48] & ~x[51] & ~x[54] & ~x[55] & ~x[59];
			partial_clause[26] 	= partial_clause_prev[26] & 1'b1;
			partial_clause[27] 	= partial_clause_prev[27] & ~x[15] & ~x[18] & ~x[29] & ~x[51] & ~x[52] & ~x[55];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[21] & ~x[40] & ~x[45] & ~x[49];
			partial_clause[29] 	= partial_clause_prev[29] & ~x[2] & ~x[16] & ~x[21] & ~x[22] & ~x[25] & ~x[48] & ~x[49] & ~x[57] & ~x[59] & ~x[63];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[1] & ~x[14];
			partial_clause[31] 	= partial_clause_prev[31] & ~x[21] & ~x[43] & ~x[46];
			partial_clause[32] 	= partial_clause_prev[32] & ~x[2] & ~x[9] & ~x[22] & ~x[28] & ~x[33] & ~x[34] & ~x[44] & ~x[56] & ~x[63];
			partial_clause[33] 	= partial_clause_prev[33] & 1'b1;
			partial_clause[34] 	= partial_clause_prev[34] & ~x[13] & ~x[16] & ~x[18] & ~x[25] & ~x[29] & ~x[35] & ~x[36] & ~x[37] & ~x[40] & ~x[42] & ~x[44] & ~x[49] & ~x[52] & ~x[53];
			partial_clause[35] 	= partial_clause_prev[35] & ~x[4] & ~x[21] & ~x[24] & ~x[32] & ~x[54] & ~x[56];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[6] & ~x[10] & ~x[12] & ~x[21] & ~x[34] & ~x[41] & ~x[42] & ~x[54];
			partial_clause[37] 	= partial_clause_prev[37] & ~x[6] & ~x[23] & ~x[25] & ~x[33] & ~x[48];
			partial_clause[38] 	= partial_clause_prev[38] & ~x[5] & ~x[24] & ~x[29] & ~x[52] & ~x[55] & ~x[57];
			partial_clause[39] 	= partial_clause_prev[39] & ~x[24] & ~x[32] & ~x[35];
			partial_clause[40] 	= partial_clause_prev[40] & ~x[2] & ~x[9] & ~x[26] & ~x[52];
			partial_clause[41] 	= partial_clause_prev[41] & 1'b1;
			partial_clause[42] 	= partial_clause_prev[42] & ~x[10] & ~x[14] & ~x[27];
			partial_clause[43] 	= partial_clause_prev[43] & ~x[10] & ~x[18] & ~x[34];
			partial_clause[44] 	= partial_clause_prev[44] & ~x[5] & ~x[41] & ~x[45];
			partial_clause[45] 	= partial_clause_prev[45] & ~x[9];
			partial_clause[46] 	= partial_clause_prev[46] & ~x[7] & ~x[14] & ~x[16] & ~x[20] & ~x[25] & ~x[30] & ~x[42] & ~x[44] & ~x[47] & ~x[51] & ~x[63];
			partial_clause[47] 	= partial_clause_prev[47] & ~x[7] & ~x[16] & ~x[32] & ~x[35] & ~x[52] & ~x[53] & ~x[61];
			partial_clause[48] 	= partial_clause_prev[48] & x[60];
			partial_clause[49] 	= partial_clause_prev[49] & 1'b1;
			partial_clause[50] 	= partial_clause_prev[50] & ~x[0] & ~x[11];
			partial_clause[51] 	= partial_clause_prev[51] & 1'b1;
			partial_clause[52] 	= partial_clause_prev[52] & 1'b1;
			partial_clause[53] 	= partial_clause_prev[53] & 1'b1;
			partial_clause[54] 	= partial_clause_prev[54] & ~x[63];
			partial_clause[55] 	= partial_clause_prev[55] & 1'b1;
			partial_clause[56] 	= partial_clause_prev[56] & 1'b1;
			partial_clause[57] 	= partial_clause_prev[57] & ~x[13] & ~x[23] & ~x[24] & ~x[26] & ~x[28] & ~x[29] & ~x[30] & ~x[38] & ~x[40] & ~x[44] & ~x[51] & ~x[53] & ~x[54] & ~x[55];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[0] & ~x[5] & ~x[6] & ~x[20] & ~x[48];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[1] & ~x[2] & ~x[11] & ~x[19] & ~x[24] & ~x[29] & ~x[30] & ~x[39] & ~x[41] & ~x[49] & ~x[53] & ~x[56] & ~x[60] & ~x[63];
			partial_clause[60] 	= partial_clause_prev[60] & 1'b1;
			partial_clause[61] 	= partial_clause_prev[61] & ~x[55];
			partial_clause[62] 	= partial_clause_prev[62] & ~x[6] & ~x[26] & ~x[30] & ~x[44] & ~x[46];
			partial_clause[63] 	= partial_clause_prev[63] & ~x[8] & ~x[45];
			partial_clause[64] 	= partial_clause_prev[64] & ~x[61];
			partial_clause[65] 	= partial_clause_prev[65] & ~x[11];
			partial_clause[66] 	= partial_clause_prev[66] & 1'b1;
			partial_clause[67] 	= partial_clause_prev[67] & 1'b1;
			partial_clause[68] 	= partial_clause_prev[68] & 1'b1;
			partial_clause[69] 	= partial_clause_prev[69] & ~x[3] & ~x[12] & ~x[23] & ~x[24] & ~x[35] & ~x[36] & ~x[42] & ~x[45] & ~x[48] & ~x[52] & ~x[53];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[4] & ~x[12] & ~x[13] & ~x[18] & ~x[27] & ~x[31] & ~x[34] & ~x[39] & ~x[59];
			partial_clause[71] 	= partial_clause_prev[71] & ~x[14] & ~x[18] & ~x[21] & ~x[27];
			partial_clause[72] 	= partial_clause_prev[72] & ~x[43];
			partial_clause[73] 	= partial_clause_prev[73] & ~x[34];
			partial_clause[74] 	= partial_clause_prev[74] & ~x[1] & ~x[3] & ~x[6] & ~x[9] & ~x[11] & ~x[12] & ~x[24] & ~x[31];
			partial_clause[75] 	= partial_clause_prev[75] & ~x[5];
			partial_clause[76] 	= partial_clause_prev[76] & ~x[2] & ~x[4] & ~x[12] & ~x[13] & ~x[14] & ~x[16] & ~x[17] & ~x[26] & ~x[28] & ~x[35] & ~x[39] & ~x[42] & ~x[44] & ~x[48] & ~x[49] & ~x[53];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[26];
			partial_clause[78] 	= partial_clause_prev[78] & ~x[12];
			partial_clause[79] 	= partial_clause_prev[79] & ~x[8] & ~x[14] & ~x[15] & ~x[19] & ~x[28] & ~x[35] & ~x[42] & ~x[46] & ~x[47] & ~x[62];
			partial_clause[80] 	= partial_clause_prev[80] & 1'b1;
			partial_clause[81] 	= partial_clause_prev[81] & ~x[3] & ~x[28] & ~x[54];
			partial_clause[82] 	= partial_clause_prev[82] & 1'b1;
			partial_clause[83] 	= partial_clause_prev[83] & 1'b1;
			partial_clause[84] 	= partial_clause_prev[84] & ~x[14] & ~x[22] & ~x[27] & ~x[29];
			partial_clause[85] 	= partial_clause_prev[85] & ~x[14] & ~x[15] & ~x[17] & ~x[22] & ~x[27] & ~x[28] & ~x[35] & ~x[36] & ~x[48] & ~x[56] & ~x[59] & ~x[60] & ~x[63];
			partial_clause[86] 	= partial_clause_prev[86] & ~x[5] & ~x[12] & ~x[22] & ~x[25] & ~x[32] & ~x[42] & ~x[55];
			partial_clause[87] 	= partial_clause_prev[87] & ~x[0] & ~x[4] & ~x[10] & ~x[13] & ~x[21] & ~x[26] & ~x[40] & ~x[53];
			partial_clause[88] 	= partial_clause_prev[88] & ~x[1] & ~x[5] & ~x[14] & ~x[20] & ~x[23] & ~x[26] & ~x[28] & ~x[38] & ~x[39] & ~x[40] & ~x[42] & ~x[49] & ~x[50] & ~x[56];
			partial_clause[89] 	= partial_clause_prev[89] & ~x[7] & ~x[12] & ~x[15] & ~x[45] & ~x[51];
			partial_clause[90] 	= partial_clause_prev[90] & 1'b1;
			partial_clause[91] 	= partial_clause_prev[91] & ~x[10] & ~x[23] & ~x[26];
			partial_clause[92] 	= partial_clause_prev[92] & ~x[49] & ~x[54];
			partial_clause[93] 	= partial_clause_prev[93] & ~x[2] & ~x[3] & ~x[5] & ~x[7] & ~x[13] & ~x[16] & ~x[22] & ~x[23] & ~x[27] & ~x[28] & ~x[29] & ~x[44] & ~x[47] & ~x[50] & ~x[55];
			partial_clause[94] 	= partial_clause_prev[94] & 1'b1;
			partial_clause[95] 	= partial_clause_prev[95] & ~x[5] & ~x[7] & ~x[9] & ~x[16] & ~x[18] & ~x[21] & ~x[23] & ~x[24] & ~x[25] & ~x[26] & ~x[32] & ~x[33] & ~x[35] & ~x[36] & ~x[37] & ~x[42] & ~x[43] & ~x[45] & ~x[59];
			partial_clause[96] 	= partial_clause_prev[96] & 1'b1;
			partial_clause[97] 	= partial_clause_prev[97] & ~x[6] & ~x[10] & ~x[11] & ~x[13] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[20] & ~x[28] & ~x[29] & ~x[36] & ~x[40] & ~x[41] & ~x[42] & ~x[44] & ~x[50];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[3] & ~x[4] & ~x[7] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[26] & ~x[27] & ~x[31] & ~x[33] & ~x[37] & ~x[40] & ~x[50] & ~x[56];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[0] & ~x[6] & ~x[7] & ~x[10] & ~x[14] & ~x[17] & ~x[18] & ~x[23] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & ~x[30] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[41] & ~x[42] & ~x[44] & ~x[45] & ~x[46] & ~x[48] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[100] 	= partial_clause_prev[100] & ~x[0];
			partial_clause[101] 	= partial_clause_prev[101] & 1'b1;
			partial_clause[102] 	= partial_clause_prev[102] & ~x[29] & ~x[56];
			partial_clause[103] 	= partial_clause_prev[103] & ~x[2] & ~x[6] & ~x[10] & ~x[12] & ~x[14] & ~x[15] & ~x[17] & ~x[20] & ~x[21] & ~x[23] & ~x[26] & ~x[27] & ~x[31] & ~x[33] & ~x[34] & ~x[47] & ~x[48] & ~x[49] & ~x[52] & ~x[53] & ~x[55] & ~x[57] & ~x[58];
			partial_clause[104] 	= partial_clause_prev[104] & ~x[9] & ~x[12] & ~x[15] & ~x[39] & ~x[43] & ~x[53] & ~x[55] & ~x[57] & ~x[62] & ~x[63];
			partial_clause[105] 	= partial_clause_prev[105] & ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[7] & ~x[9] & ~x[16] & ~x[17] & ~x[25] & ~x[33] & ~x[39] & ~x[40] & ~x[46] & ~x[47] & ~x[50] & ~x[55] & ~x[62];
			partial_clause[106] 	= partial_clause_prev[106] & ~x[3] & ~x[16] & ~x[40] & ~x[46] & ~x[47] & ~x[53] & ~x[58];
			partial_clause[107] 	= partial_clause_prev[107] & ~x[5] & ~x[6] & ~x[10] & ~x[14] & ~x[18] & ~x[30] & ~x[34] & ~x[35] & ~x[44] & ~x[46] & ~x[49] & ~x[63];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[0] & ~x[5] & ~x[9] & ~x[11] & ~x[18] & ~x[19] & ~x[24] & ~x[32] & ~x[33] & ~x[48] & ~x[51] & ~x[52] & ~x[53] & ~x[56] & ~x[57];
			partial_clause[109] 	= partial_clause_prev[109] & ~x[63];
			partial_clause[110] 	= partial_clause_prev[110] & ~x[54];
			partial_clause[111] 	= partial_clause_prev[111] & 1'b1;
			partial_clause[112] 	= partial_clause_prev[112] & ~x[40] & ~x[48];
			partial_clause[113] 	= partial_clause_prev[113] & ~x[59];
			partial_clause[114] 	= partial_clause_prev[114] & 1'b1;
			partial_clause[115] 	= partial_clause_prev[115] & ~x[2] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[12] & ~x[13] & ~x[14] & ~x[17] & ~x[19] & ~x[33] & ~x[35] & ~x[36] & ~x[37] & ~x[46] & ~x[50] & ~x[51] & ~x[56];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[1] & ~x[15] & ~x[22] & ~x[24] & ~x[32] & ~x[34] & ~x[35] & ~x[40] & ~x[46] & ~x[50] & ~x[58];
			partial_clause[117] 	= partial_clause_prev[117] & 1'b1;
			partial_clause[118] 	= partial_clause_prev[118] & ~x[13] & ~x[32] & ~x[35] & ~x[36] & ~x[41] & ~x[43] & ~x[44] & ~x[47] & ~x[51] & ~x[59];
			partial_clause[119] 	= partial_clause_prev[119] & ~x[1] & ~x[4] & ~x[12] & ~x[23] & ~x[24] & ~x[28] & ~x[29] & ~x[32] & ~x[35] & ~x[36] & ~x[49] & ~x[51] & ~x[63];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[0] & ~x[1] & ~x[2] & ~x[4] & ~x[6] & ~x[9] & ~x[10] & ~x[12] & ~x[14] & ~x[15] & ~x[17] & ~x[22] & ~x[23] & ~x[28] & ~x[29] & ~x[30] & ~x[34] & ~x[37] & ~x[39] & ~x[40] & ~x[41] & ~x[43] & ~x[47] & ~x[49] & ~x[52] & ~x[53] & ~x[54] & ~x[55];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[12] & ~x[14] & ~x[17] & ~x[24] & ~x[44] & ~x[47] & ~x[49] & ~x[52];
			partial_clause[122] 	= partial_clause_prev[122] & ~x[11] & ~x[16] & ~x[30] & ~x[44] & ~x[46] & ~x[60];
			partial_clause[123] 	= partial_clause_prev[123] & ~x[0] & ~x[2] & ~x[15] & ~x[18] & ~x[22] & ~x[29] & ~x[32] & ~x[41] & ~x[47] & ~x[49] & ~x[56] & ~x[58];
			partial_clause[124] 	= partial_clause_prev[124] & 1'b1;
			partial_clause[125] 	= partial_clause_prev[125] & ~x[39] & ~x[45];
			partial_clause[126] 	= partial_clause_prev[126] & ~x[7] & ~x[31] & ~x[32] & ~x[40] & ~x[56] & ~x[58] & ~x[61];
			partial_clause[127] 	= partial_clause_prev[127] & ~x[2] & ~x[7] & ~x[8] & ~x[13] & ~x[14] & ~x[17] & ~x[18] & ~x[20] & ~x[21] & ~x[24] & ~x[25] & ~x[27] & ~x[28] & ~x[30] & ~x[35] & ~x[37] & ~x[38] & ~x[41] & ~x[43] & ~x[44] & ~x[45] & ~x[52] & ~x[56] & ~x[62];
			partial_clause[128] 	= partial_clause_prev[128] & ~x[20] & ~x[28] & ~x[29] & ~x[31] & ~x[34] & ~x[53] & ~x[60] & ~x[62];
			partial_clause[129] 	= partial_clause_prev[129] & ~x[2] & ~x[8] & ~x[11] & ~x[14] & ~x[16] & ~x[21] & ~x[31] & ~x[32] & ~x[34] & ~x[35] & ~x[42] & ~x[43] & ~x[44] & ~x[52] & ~x[56] & ~x[62];
			partial_clause[130] 	= partial_clause_prev[130] & ~x[2] & ~x[8] & ~x[10] & ~x[14] & ~x[16] & ~x[41] & ~x[47] & ~x[49] & ~x[52] & ~x[56];
			partial_clause[131] 	= partial_clause_prev[131] & ~x[25];
			partial_clause[132] 	= partial_clause_prev[132] & ~x[7] & ~x[19] & ~x[25] & ~x[40] & ~x[46];
			partial_clause[133] 	= partial_clause_prev[133] & ~x[50];
			partial_clause[134] 	= partial_clause_prev[134] & ~x[0] & ~x[1] & ~x[4] & ~x[9] & ~x[15] & ~x[17] & ~x[18] & ~x[19] & ~x[25] & ~x[28] & ~x[35] & ~x[40] & ~x[41] & ~x[44] & ~x[45] & ~x[47] & ~x[50] & ~x[55] & ~x[56];
			partial_clause[135] 	= partial_clause_prev[135] & ~x[22] & ~x[27] & ~x[41] & ~x[46] & ~x[53];
			partial_clause[136] 	= partial_clause_prev[136] & ~x[3] & ~x[5] & ~x[12] & ~x[17] & ~x[20] & ~x[30] & ~x[37] & ~x[38] & ~x[41] & ~x[42] & ~x[47] & ~x[51] & ~x[55];
			partial_clause[137] 	= partial_clause_prev[137] & ~x[30] & ~x[63];
			partial_clause[138] 	= partial_clause_prev[138] & ~x[38] & ~x[44];
			partial_clause[139] 	= partial_clause_prev[139] & ~x[1] & ~x[3] & ~x[5] & ~x[9] & ~x[10] & ~x[22] & ~x[24] & ~x[25] & ~x[29] & ~x[33] & ~x[35] & ~x[45] & ~x[46] & ~x[47];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[9] & ~x[10] & ~x[14] & ~x[15] & ~x[16] & ~x[24] & ~x[27] & ~x[43] & ~x[45] & ~x[46] & ~x[51] & ~x[53] & ~x[56];
			partial_clause[141] 	= partial_clause_prev[141] & ~x[3] & ~x[26] & ~x[32] & ~x[43] & ~x[44] & ~x[49] & ~x[51] & ~x[55];
			partial_clause[142] 	= partial_clause_prev[142] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[19] & ~x[27] & ~x[29] & ~x[32] & ~x[40] & ~x[42] & ~x[47] & ~x[62];
			partial_clause[143] 	= partial_clause_prev[143] & ~x[14] & ~x[20] & ~x[22] & ~x[53];
			partial_clause[144] 	= partial_clause_prev[144] & ~x[0] & ~x[9] & ~x[10] & ~x[13] & ~x[14] & ~x[15] & ~x[22] & ~x[30] & ~x[44] & ~x[48];
			partial_clause[145] 	= partial_clause_prev[145] & ~x[34];
			partial_clause[146] 	= partial_clause_prev[146] & ~x[10] & ~x[17] & ~x[20] & ~x[23] & ~x[27] & ~x[28] & ~x[31] & ~x[37] & ~x[43] & ~x[44] & ~x[58];
			partial_clause[147] 	= partial_clause_prev[147] & ~x[14] & ~x[22] & ~x[27] & ~x[42] & ~x[47] & ~x[49] & ~x[51] & ~x[52];
			partial_clause[148] 	= partial_clause_prev[148] & ~x[4] & ~x[12] & ~x[18] & ~x[27] & ~x[32] & ~x[39] & ~x[42] & ~x[43] & ~x[45] & ~x[56] & ~x[58];
			partial_clause[149] 	= partial_clause_prev[149] & ~x[30] & ~x[37];
			partial_clause[150] 	= partial_clause_prev[150] & ~x[10] & ~x[18] & ~x[30] & ~x[36] & ~x[56];
			partial_clause[151] 	= partial_clause_prev[151] & ~x[15];
			partial_clause[152] 	= partial_clause_prev[152] & ~x[6] & ~x[10] & ~x[12] & ~x[27] & ~x[29] & ~x[31] & ~x[34] & ~x[42];
			partial_clause[153] 	= partial_clause_prev[153] & ~x[2] & ~x[13] & ~x[26] & ~x[45] & ~x[47] & ~x[49];
			partial_clause[154] 	= partial_clause_prev[154] & ~x[60];
			partial_clause[155] 	= partial_clause_prev[155] & 1'b1;
			partial_clause[156] 	= partial_clause_prev[156] & 1'b1;
			partial_clause[157] 	= partial_clause_prev[157] & 1'b1;
			partial_clause[158] 	= partial_clause_prev[158] & ~x[0] & ~x[6] & ~x[7] & ~x[10] & ~x[16] & ~x[19] & ~x[20] & ~x[23] & ~x[24] & ~x[26] & ~x[32] & ~x[34] & ~x[39] & ~x[41] & ~x[44] & ~x[45] & ~x[47] & ~x[61] & ~x[62];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[12] & ~x[13] & ~x[31] & ~x[32] & ~x[40] & ~x[41] & ~x[46] & ~x[50] & ~x[53];
			partial_clause[160] 	= partial_clause_prev[160] & ~x[1] & ~x[9] & ~x[10] & ~x[26] & ~x[35] & ~x[59];
			partial_clause[161] 	= partial_clause_prev[161] & ~x[0] & ~x[9] & ~x[12] & ~x[18] & ~x[19] & ~x[28] & ~x[36] & ~x[38] & ~x[57];
			partial_clause[162] 	= partial_clause_prev[162] & ~x[9] & ~x[20] & ~x[23] & ~x[25] & ~x[45] & ~x[63];
			partial_clause[163] 	= partial_clause_prev[163] & ~x[5];
			partial_clause[164] 	= partial_clause_prev[164] & ~x[28] & ~x[29] & ~x[36] & ~x[37];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[10] & ~x[20] & ~x[30] & ~x[35] & ~x[37] & ~x[42] & ~x[57];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[1] & ~x[3] & ~x[6] & ~x[24] & ~x[27] & ~x[29] & ~x[31] & ~x[38] & ~x[40] & ~x[51] & ~x[52];
			partial_clause[167] 	= partial_clause_prev[167] & ~x[52];
			partial_clause[168] 	= partial_clause_prev[168] & 1'b1;
			partial_clause[169] 	= partial_clause_prev[169] & 1'b1;
			partial_clause[170] 	= partial_clause_prev[170] & 1'b1;
			partial_clause[171] 	= partial_clause_prev[171] & ~x[1] & ~x[7] & ~x[11] & ~x[30] & ~x[41] & ~x[59];
			partial_clause[172] 	= partial_clause_prev[172] & ~x[34];
			partial_clause[173] 	= partial_clause_prev[173] & ~x[6] & ~x[17] & ~x[20] & ~x[21] & ~x[26] & ~x[27] & ~x[29] & ~x[31] & ~x[59];
			partial_clause[174] 	= partial_clause_prev[174] & ~x[7] & ~x[34] & ~x[60];
			partial_clause[175] 	= partial_clause_prev[175] & ~x[62] & ~x[63];
			partial_clause[176] 	= partial_clause_prev[176] & 1'b1;
			partial_clause[177] 	= partial_clause_prev[177] & ~x[9] & ~x[17] & ~x[32] & ~x[40] & ~x[53];
			partial_clause[178] 	= partial_clause_prev[178] & ~x[0] & ~x[16] & ~x[21] & ~x[39];
			partial_clause[179] 	= partial_clause_prev[179] & 1'b1;
			partial_clause[180] 	= partial_clause_prev[180] & ~x[9] & ~x[50];
			partial_clause[181] 	= partial_clause_prev[181] & 1'b1;
			partial_clause[182] 	= partial_clause_prev[182] & 1'b1;
			partial_clause[183] 	= partial_clause_prev[183] & ~x[0] & ~x[1] & ~x[14] & ~x[15] & ~x[18] & ~x[24] & ~x[35] & ~x[38] & ~x[41] & ~x[45] & ~x[47] & ~x[52] & ~x[53] & ~x[55] & ~x[56] & ~x[57] & ~x[59];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[10] & ~x[12] & ~x[13] & ~x[19] & ~x[24] & ~x[33] & ~x[38] & ~x[53] & ~x[57] & ~x[58];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[0] & ~x[18] & ~x[19] & ~x[21] & ~x[51] & ~x[52];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[10] & ~x[11] & ~x[17] & ~x[18] & ~x[24] & ~x[31] & ~x[32] & ~x[33] & ~x[36] & ~x[41] & ~x[43] & ~x[44] & ~x[45] & ~x[46] & ~x[47] & ~x[48] & ~x[59] & ~x[61] & ~x[63];
			partial_clause[187] 	= partial_clause_prev[187] & ~x[2] & ~x[7] & ~x[18] & ~x[21] & ~x[33] & ~x[36] & ~x[39] & ~x[44] & ~x[46] & ~x[48];
			partial_clause[188] 	= partial_clause_prev[188] & 1'b1;
			partial_clause[189] 	= partial_clause_prev[189] & 1'b1;
			partial_clause[190] 	= partial_clause_prev[190] & ~x[10] & ~x[29] & ~x[35] & ~x[40];
			partial_clause[191] 	= partial_clause_prev[191] & ~x[52] & ~x[58] & ~x[61];
			partial_clause[192] 	= partial_clause_prev[192] & ~x[2] & ~x[8] & ~x[10] & ~x[21] & ~x[33] & ~x[42];
			partial_clause[193] 	= partial_clause_prev[193] & ~x[0] & ~x[17] & ~x[26] & ~x[36] & ~x[52] & ~x[53];
			partial_clause[194] 	= partial_clause_prev[194] & ~x[20] & ~x[54] & ~x[58];
			partial_clause[195] 	= partial_clause_prev[195] & ~x[2] & ~x[3] & ~x[6] & ~x[12] & ~x[13] & ~x[14] & ~x[18] & ~x[30] & ~x[34] & ~x[36] & ~x[53] & ~x[56] & ~x[58];
			partial_clause[196] 	= partial_clause_prev[196] & ~x[48];
			partial_clause[197] 	= partial_clause_prev[197] & ~x[4] & ~x[12] & ~x[14] & ~x[17] & ~x[18] & ~x[35] & ~x[38] & ~x[41] & ~x[42] & ~x[52] & ~x[59];
			partial_clause[198] 	= partial_clause_prev[198] & 1'b1;
			partial_clause[199] 	= partial_clause_prev[199] & 1'b1;
			partial_clause[200] 	= partial_clause_prev[200] & ~x[24] & ~x[27] & ~x[35] & ~x[46];
			partial_clause[201] 	= partial_clause_prev[201] & ~x[11] & ~x[22] & ~x[23] & ~x[31] & ~x[37] & ~x[39] & ~x[44] & ~x[46] & ~x[53] & ~x[59] & ~x[62] & ~x[63];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[0] & ~x[1] & ~x[2] & ~x[4] & ~x[16] & ~x[18] & ~x[25] & ~x[31] & ~x[32] & ~x[42] & ~x[44] & ~x[45] & ~x[49];
			partial_clause[203] 	= partial_clause_prev[203] & ~x[47];
			partial_clause[204] 	= partial_clause_prev[204] & ~x[0] & ~x[5] & ~x[7] & ~x[12] & ~x[18] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[28] & ~x[29] & ~x[39] & ~x[41] & ~x[44] & ~x[56] & ~x[58];
			partial_clause[205] 	= partial_clause_prev[205] & ~x[10];
			partial_clause[206] 	= partial_clause_prev[206] & ~x[0] & ~x[2] & ~x[4] & ~x[6] & ~x[9] & ~x[14] & ~x[15] & ~x[18] & ~x[19] & ~x[21] & ~x[23] & ~x[28] & ~x[29] & ~x[37] & ~x[41] & ~x[50] & ~x[53] & ~x[54] & ~x[56];
			partial_clause[207] 	= partial_clause_prev[207] & ~x[4] & ~x[9] & ~x[11] & ~x[19] & ~x[26] & ~x[39] & ~x[46] & ~x[47] & ~x[53] & ~x[54];
			partial_clause[208] 	= partial_clause_prev[208] & ~x[1] & ~x[8] & ~x[9] & ~x[14] & ~x[22] & ~x[32] & ~x[52] & ~x[56] & ~x[58];
			partial_clause[209] 	= partial_clause_prev[209] & 1'b1;
			partial_clause[210] 	= partial_clause_prev[210] & ~x[2] & ~x[10] & ~x[19] & ~x[22] & ~x[25] & ~x[40] & ~x[43] & ~x[44] & ~x[55] & ~x[56];
			partial_clause[211] 	= partial_clause_prev[211] & 1'b1;
			partial_clause[212] 	= partial_clause_prev[212] & ~x[43] & ~x[54];
			partial_clause[213] 	= partial_clause_prev[213] & 1'b1;
			partial_clause[214] 	= partial_clause_prev[214] & ~x[16];
			partial_clause[215] 	= partial_clause_prev[215] & 1'b1;
			partial_clause[216] 	= partial_clause_prev[216] & ~x[1] & ~x[3] & ~x[16] & ~x[17];
			partial_clause[217] 	= partial_clause_prev[217] & ~x[2] & ~x[19] & ~x[24] & ~x[27] & ~x[28] & ~x[45] & ~x[51];
			partial_clause[218] 	= partial_clause_prev[218] & ~x[58];
			partial_clause[219] 	= partial_clause_prev[219] & ~x[50] & ~x[51];
			partial_clause[220] 	= partial_clause_prev[220] & ~x[0] & ~x[2] & ~x[4] & ~x[7] & ~x[9] & ~x[13] & ~x[15] & ~x[20] & ~x[21] & ~x[24] & ~x[27] & ~x[30] & ~x[33] & ~x[35] & ~x[42] & ~x[43] & ~x[45];
			partial_clause[221] 	= partial_clause_prev[221] & ~x[16] & ~x[47];
			partial_clause[222] 	= partial_clause_prev[222] & ~x[16];
			partial_clause[223] 	= partial_clause_prev[223] & ~x[21] & ~x[42];
			partial_clause[224] 	= partial_clause_prev[224] & ~x[5] & ~x[7] & ~x[34] & ~x[36] & ~x[48] & ~x[58] & ~x[59];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[42] & ~x[47];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[8] & ~x[10] & ~x[11] & ~x[12] & ~x[14] & ~x[16] & ~x[17] & ~x[20] & ~x[23] & ~x[26] & ~x[28] & ~x[29] & ~x[30] & ~x[31] & ~x[32] & ~x[39] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[47] & ~x[49] & ~x[51] & ~x[53] & ~x[58] & ~x[61];
			partial_clause[227] 	= partial_clause_prev[227] & 1'b1;
			partial_clause[228] 	= partial_clause_prev[228] & ~x[5] & ~x[7] & ~x[9] & ~x[10] & ~x[22] & ~x[29] & ~x[33] & ~x[36] & ~x[39] & ~x[40] & ~x[42] & ~x[52] & ~x[57];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[3] & ~x[15] & ~x[19] & ~x[26] & ~x[28] & ~x[29] & ~x[30] & ~x[46] & ~x[51] & ~x[53] & ~x[56] & ~x[58];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[0] & ~x[4] & ~x[5] & ~x[6] & ~x[13] & ~x[14] & ~x[16] & ~x[19] & ~x[20] & ~x[23] & ~x[24] & ~x[27] & ~x[28] & ~x[30] & ~x[31] & ~x[33] & ~x[41] & ~x[44] & ~x[46] & ~x[50] & ~x[52] & ~x[58] & ~x[59];
			partial_clause[231] 	= partial_clause_prev[231] & ~x[19] & ~x[21] & ~x[29] & ~x[46];
			partial_clause[232] 	= partial_clause_prev[232] & 1'b1;
			partial_clause[233] 	= partial_clause_prev[233] & ~x[55];
			partial_clause[234] 	= partial_clause_prev[234] & ~x[37];
			partial_clause[235] 	= partial_clause_prev[235] & 1'b1;
			partial_clause[236] 	= partial_clause_prev[236] & 1'b1;
			partial_clause[237] 	= partial_clause_prev[237] & 1'b1;
			partial_clause[238] 	= partial_clause_prev[238] & ~x[41] & ~x[58];
			partial_clause[239] 	= partial_clause_prev[239] & ~x[21] & ~x[22] & ~x[24] & ~x[38];
			partial_clause[240] 	= partial_clause_prev[240] & ~x[2] & ~x[12] & ~x[17] & ~x[20] & ~x[34] & ~x[36] & ~x[40] & ~x[63];
			partial_clause[241] 	= partial_clause_prev[241] & ~x[2] & ~x[14] & ~x[37] & ~x[38] & ~x[41];
			partial_clause[242] 	= partial_clause_prev[242] & ~x[1] & ~x[4] & ~x[8] & ~x[9] & ~x[10] & ~x[16] & ~x[20] & ~x[22] & ~x[25] & ~x[38] & ~x[51] & ~x[53] & ~x[63];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[14] & ~x[19] & ~x[23] & ~x[26] & ~x[37] & ~x[39] & ~x[46] & ~x[54];
			partial_clause[244] 	= partial_clause_prev[244] & ~x[18] & ~x[51] & ~x[53] & ~x[57];
			partial_clause[245] 	= partial_clause_prev[245] & 1'b1;
			partial_clause[246] 	= partial_clause_prev[246] & ~x[6] & ~x[10] & ~x[31] & ~x[50];
			partial_clause[247] 	= partial_clause_prev[247] & ~x[0] & ~x[1] & ~x[4] & ~x[10] & ~x[11] & ~x[14] & ~x[15] & ~x[22] & ~x[23] & ~x[25] & ~x[31] & ~x[32] & ~x[37] & ~x[42] & ~x[45] & ~x[48] & ~x[50] & ~x[51] & ~x[53] & ~x[56] & ~x[61] & ~x[62];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[1] & ~x[2] & ~x[4] & ~x[11] & ~x[12] & ~x[13] & ~x[17] & ~x[18] & ~x[19] & ~x[28] & ~x[29] & ~x[30] & ~x[38] & ~x[39] & ~x[41] & ~x[42] & ~x[43] & ~x[47] & ~x[50] & ~x[53] & ~x[54] & ~x[55];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[16] & ~x[43];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[0] & ~x[3] & ~x[5] & ~x[7] & ~x[9] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[23] & ~x[24] & ~x[25] & ~x[27] & ~x[28] & ~x[30] & ~x[31] & ~x[33] & ~x[34] & ~x[36] & ~x[37] & ~x[40] & ~x[45] & ~x[46] & ~x[47] & ~x[50] & ~x[53] & ~x[55] & ~x[56] & ~x[59] & ~x[60] & ~x[61];
			partial_clause[251] 	= partial_clause_prev[251] & ~x[36];
			partial_clause[252] 	= partial_clause_prev[252] & ~x[1] & ~x[2] & ~x[5] & ~x[8] & ~x[9] & ~x[11] & ~x[12] & ~x[14] & ~x[17] & ~x[19] & ~x[22] & ~x[45] & ~x[50] & ~x[54];
			partial_clause[253] 	= partial_clause_prev[253] & ~x[10] & ~x[22] & ~x[24] & ~x[38] & ~x[49];
			partial_clause[254] 	= partial_clause_prev[254] & ~x[0] & ~x[23] & ~x[27] & ~x[37] & ~x[44] & ~x[51] & ~x[52];
			partial_clause[255] 	= partial_clause_prev[255] & ~x[19] & ~x[21] & ~x[49];
			partial_clause[256] 	= partial_clause_prev[256] & 1'b1;
			partial_clause[257] 	= partial_clause_prev[257] & ~x[4] & ~x[10] & ~x[17] & ~x[28] & ~x[31] & ~x[32] & ~x[33] & ~x[43] & ~x[63];
			partial_clause[258] 	= partial_clause_prev[258] & ~x[8] & ~x[16] & ~x[21] & ~x[23] & ~x[24] & ~x[26] & ~x[33] & ~x[35] & ~x[41] & ~x[51] & ~x[57] & ~x[63];
			partial_clause[259] 	= partial_clause_prev[259] & 1'b1;
			partial_clause[260] 	= partial_clause_prev[260] & ~x[5] & ~x[20] & ~x[29] & ~x[30] & ~x[44] & ~x[55];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[18] & ~x[30] & ~x[31] & ~x[35] & ~x[43] & ~x[49] & ~x[53] & ~x[57];
			partial_clause[262] 	= partial_clause_prev[262] & ~x[22] & ~x[53];
			partial_clause[263] 	= partial_clause_prev[263] & ~x[0] & ~x[22] & ~x[49] & ~x[61];
			partial_clause[264] 	= partial_clause_prev[264] & ~x[56];
			partial_clause[265] 	= partial_clause_prev[265] & 1'b1;
			partial_clause[266] 	= partial_clause_prev[266] & ~x[6] & ~x[9] & ~x[10] & ~x[16] & ~x[18] & ~x[24] & ~x[27] & ~x[32] & ~x[33] & ~x[38] & ~x[40] & ~x[53] & ~x[54] & ~x[55] & ~x[59];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[0] & ~x[1] & ~x[5] & ~x[6] & ~x[12] & ~x[16] & ~x[21] & ~x[24] & ~x[27] & ~x[32] & ~x[33] & ~x[36] & ~x[37] & ~x[42] & ~x[44] & ~x[50] & ~x[52] & ~x[54] & ~x[55] & ~x[58] & ~x[60];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[0] & ~x[3] & ~x[6] & ~x[7] & ~x[10] & ~x[11] & ~x[14] & ~x[17] & ~x[19] & ~x[26] & ~x[30] & ~x[34] & ~x[37] & ~x[38] & ~x[39] & ~x[41] & ~x[42] & ~x[47] & ~x[50] & ~x[52] & ~x[54] & ~x[56] & ~x[57] & ~x[58] & ~x[60];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[1] & ~x[2] & ~x[7] & ~x[8] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[21] & ~x[25] & ~x[27] & ~x[28] & ~x[31] & ~x[41] & ~x[46] & ~x[48] & ~x[52] & ~x[53] & ~x[55] & ~x[57] & ~x[59];
			partial_clause[270] 	= partial_clause_prev[270] & 1'b1;
			partial_clause[271] 	= partial_clause_prev[271] & 1'b1;
			partial_clause[272] 	= partial_clause_prev[272] & ~x[0] & ~x[6] & ~x[9] & ~x[25] & ~x[27] & ~x[28] & ~x[31] & ~x[33] & ~x[41] & ~x[50];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[3] & ~x[6] & ~x[7] & ~x[13] & ~x[14] & ~x[16] & ~x[17] & ~x[18] & ~x[20] & ~x[21] & ~x[24] & ~x[27] & ~x[29] & ~x[30] & ~x[34] & ~x[41] & ~x[48] & ~x[51] & ~x[53] & ~x[57] & ~x[58] & ~x[60];
			partial_clause[274] 	= partial_clause_prev[274] & ~x[6] & ~x[7] & ~x[14] & ~x[20] & ~x[40] & ~x[42] & ~x[44] & ~x[47] & ~x[49];
			partial_clause[275] 	= partial_clause_prev[275] & ~x[35];
			partial_clause[276] 	= partial_clause_prev[276] & ~x[1] & ~x[8] & ~x[16] & ~x[18] & ~x[24] & ~x[25] & ~x[40];
			partial_clause[277] 	= partial_clause_prev[277] & ~x[2] & ~x[17] & ~x[25] & ~x[27] & ~x[32] & ~x[33] & ~x[46] & ~x[61] & ~x[62];
			partial_clause[278] 	= partial_clause_prev[278] & 1'b1;
			partial_clause[279] 	= partial_clause_prev[279] & ~x[2] & ~x[4] & ~x[10] & ~x[12] & ~x[13] & ~x[18] & ~x[19] & ~x[28] & ~x[30] & ~x[34] & ~x[35] & ~x[48] & ~x[53];
			partial_clause[280] 	= partial_clause_prev[280] & 1'b1;
			partial_clause[281] 	= partial_clause_prev[281] & ~x[6] & ~x[19] & ~x[29] & ~x[32] & ~x[53] & ~x[56] & ~x[58];
			partial_clause[282] 	= partial_clause_prev[282] & ~x[20];
			partial_clause[283] 	= partial_clause_prev[283] & ~x[15];
			partial_clause[284] 	= partial_clause_prev[284] & ~x[23];
			partial_clause[285] 	= partial_clause_prev[285] & 1'b1;
			partial_clause[286] 	= partial_clause_prev[286] & ~x[12] & ~x[50];
			partial_clause[287] 	= partial_clause_prev[287] & ~x[0] & ~x[1] & ~x[4] & ~x[8] & ~x[10] & ~x[15] & ~x[18] & ~x[21] & ~x[24] & ~x[25] & ~x[32] & ~x[42] & ~x[47] & ~x[56];
			partial_clause[288] 	= partial_clause_prev[288] & 1'b1;
			partial_clause[289] 	= partial_clause_prev[289] & ~x[5] & ~x[10] & ~x[35] & ~x[52];
			partial_clause[290] 	= partial_clause_prev[290] & ~x[2];
			partial_clause[291] 	= partial_clause_prev[291] & ~x[54];
			partial_clause[292] 	= partial_clause_prev[292] & ~x[10] & ~x[12] & ~x[13] & ~x[31] & ~x[35] & ~x[42] & ~x[46] & ~x[60];
			partial_clause[293] 	= partial_clause_prev[293] & ~x[27] & ~x[38] & ~x[41] & ~x[62];
			partial_clause[294] 	= partial_clause_prev[294] & ~x[30] & ~x[31] & ~x[37] & ~x[38] & ~x[55];
			partial_clause[295] 	= partial_clause_prev[295] & ~x[10] & ~x[17] & ~x[38] & ~x[39] & ~x[45];
			partial_clause[296] 	= partial_clause_prev[296] & 1'b1;
			partial_clause[297] 	= partial_clause_prev[297] & ~x[2] & ~x[3] & ~x[6] & ~x[27] & ~x[33] & ~x[39] & ~x[48] & ~x[59];
			partial_clause[298] 	= partial_clause_prev[298] & 1'b1;
			partial_clause[299] 	= partial_clause_prev[299] & ~x[29] & ~x[31] & ~x[40] & ~x[41] & ~x[51] & ~x[54];
			partial_clause[300] 	= partial_clause_prev[300] & ~x[18] & ~x[21] & ~x[24] & ~x[26] & ~x[49];
			partial_clause[301] 	= partial_clause_prev[301] & ~x[23] & ~x[24] & ~x[26] & ~x[29] & ~x[32] & ~x[35] & ~x[37] & ~x[38] & ~x[42] & ~x[45] & ~x[49] & ~x[58] & ~x[61];
			partial_clause[302] 	= partial_clause_prev[302] & ~x[27] & ~x[30] & ~x[39] & ~x[46];
			partial_clause[303] 	= partial_clause_prev[303] & ~x[8] & ~x[48] & ~x[59];
			partial_clause[304] 	= partial_clause_prev[304] & ~x[18];
			partial_clause[305] 	= partial_clause_prev[305] & ~x[18] & ~x[46] & ~x[52];
			partial_clause[306] 	= partial_clause_prev[306] & ~x[4] & ~x[35] & ~x[40] & ~x[43] & ~x[50] & ~x[61];
			partial_clause[307] 	= partial_clause_prev[307] & ~x[23] & ~x[25] & ~x[36] & ~x[43] & ~x[57];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[5] & ~x[6] & ~x[14] & ~x[15] & ~x[16] & ~x[18] & ~x[20] & ~x[30] & ~x[31] & ~x[38] & ~x[40] & ~x[44];
			partial_clause[309] 	= partial_clause_prev[309] & ~x[2] & ~x[4] & ~x[17] & ~x[23] & ~x[24] & ~x[30] & ~x[37] & ~x[38] & ~x[47] & ~x[52];
			partial_clause[310] 	= partial_clause_prev[310] & ~x[16];
			partial_clause[311] 	= partial_clause_prev[311] & ~x[31];
			partial_clause[312] 	= partial_clause_prev[312] & ~x[30];
			partial_clause[313] 	= partial_clause_prev[313] & 1'b1;
			partial_clause[314] 	= partial_clause_prev[314] & ~x[3] & ~x[37] & ~x[49];
			partial_clause[315] 	= partial_clause_prev[315] & ~x[10] & ~x[15] & ~x[26] & ~x[39] & ~x[46] & ~x[51];
			partial_clause[316] 	= partial_clause_prev[316] & ~x[1] & ~x[3] & ~x[4] & ~x[11] & ~x[14] & ~x[22] & ~x[25] & ~x[37] & ~x[51] & ~x[54];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[0] & ~x[2] & ~x[4] & ~x[15] & ~x[18] & ~x[20] & ~x[23] & ~x[51];
			partial_clause[318] 	= partial_clause_prev[318] & ~x[26] & ~x[28] & ~x[32] & ~x[33];
			partial_clause[319] 	= partial_clause_prev[319] & ~x[5] & ~x[34];
			partial_clause[320] 	= partial_clause_prev[320] & ~x[1] & ~x[3] & ~x[16] & ~x[18] & ~x[25] & ~x[26] & ~x[30] & ~x[40] & ~x[44] & ~x[45];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[8] & ~x[13] & ~x[24] & ~x[25] & ~x[27] & ~x[28] & ~x[30] & ~x[40] & ~x[45] & ~x[51];
			partial_clause[322] 	= partial_clause_prev[322] & ~x[5] & ~x[6] & ~x[7];
			partial_clause[323] 	= partial_clause_prev[323] & ~x[59];
			partial_clause[324] 	= partial_clause_prev[324] & ~x[10] & ~x[13] & ~x[31] & ~x[45];
			partial_clause[325] 	= partial_clause_prev[325] & ~x[0] & ~x[1] & ~x[4] & ~x[8] & ~x[24] & ~x[25] & ~x[27] & ~x[28] & ~x[29] & ~x[31] & ~x[43] & ~x[44] & ~x[47] & ~x[48] & ~x[50] & ~x[52] & ~x[55] & ~x[57];
			partial_clause[326] 	= partial_clause_prev[326] & ~x[3] & ~x[4] & ~x[13] & ~x[16] & ~x[24] & ~x[27] & ~x[31] & ~x[42] & ~x[43] & ~x[45] & ~x[52] & ~x[55] & ~x[57] & ~x[60] & ~x[61];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[43] & ~x[44] & ~x[47];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[2] & ~x[15] & ~x[16] & ~x[47] & ~x[51];
			partial_clause[329] 	= partial_clause_prev[329] & ~x[57];
			partial_clause[330] 	= partial_clause_prev[330] & ~x[42] & ~x[45] & ~x[46];
			partial_clause[331] 	= partial_clause_prev[331] & ~x[28] & ~x[29] & ~x[45];
			partial_clause[332] 	= partial_clause_prev[332] & ~x[4] & ~x[16] & ~x[18] & ~x[20] & ~x[38];
			partial_clause[333] 	= partial_clause_prev[333] & ~x[15] & ~x[42] & ~x[48];
			partial_clause[334] 	= partial_clause_prev[334] & ~x[2] & ~x[10] & ~x[24] & ~x[28] & ~x[29] & ~x[45] & ~x[56];
			partial_clause[335] 	= partial_clause_prev[335] & ~x[8] & ~x[9] & ~x[35] & ~x[55];
			partial_clause[336] 	= partial_clause_prev[336] & ~x[2];
			partial_clause[337] 	= partial_clause_prev[337] & ~x[0] & ~x[2] & ~x[9] & ~x[11] & ~x[15] & ~x[22] & ~x[23] & ~x[44] & ~x[46] & ~x[50];
			partial_clause[338] 	= partial_clause_prev[338] & 1'b1;
			partial_clause[339] 	= partial_clause_prev[339] & ~x[0] & ~x[2] & ~x[4] & ~x[6] & ~x[10] & ~x[13] & ~x[21] & ~x[22] & ~x[24] & ~x[25] & ~x[26] & ~x[35] & ~x[36] & ~x[37] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[45] & ~x[53] & ~x[60];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[1] & ~x[7] & ~x[14] & ~x[17] & ~x[23] & ~x[34] & ~x[39] & ~x[46] & ~x[47] & ~x[52] & ~x[54] & ~x[55] & ~x[58] & ~x[60];
			partial_clause[341] 	= partial_clause_prev[341] & 1'b1;
			partial_clause[342] 	= partial_clause_prev[342] & ~x[5] & ~x[8] & ~x[10] & ~x[13] & ~x[22] & ~x[27] & ~x[33] & ~x[34] & ~x[35] & ~x[36] & ~x[38] & ~x[49] & ~x[54] & ~x[56];
			partial_clause[343] 	= partial_clause_prev[343] & ~x[14];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[5] & ~x[9] & ~x[19] & ~x[21] & ~x[31] & ~x[48] & ~x[51] & ~x[61];
			partial_clause[345] 	= partial_clause_prev[345] & ~x[11] & ~x[26];
			partial_clause[346] 	= partial_clause_prev[346] & ~x[1] & ~x[12] & ~x[17] & ~x[30] & ~x[31] & ~x[34] & ~x[63];
			partial_clause[347] 	= partial_clause_prev[347] & ~x[1] & ~x[13] & ~x[19];
			partial_clause[348] 	= partial_clause_prev[348] & ~x[4] & ~x[12] & ~x[36];
			partial_clause[349] 	= partial_clause_prev[349] & ~x[0];
			partial_clause[350] 	= partial_clause_prev[350] & ~x[0] & ~x[3] & ~x[4] & ~x[6] & ~x[7] & ~x[9] & ~x[10] & ~x[11] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[22] & ~x[25] & ~x[27] & ~x[28] & ~x[29] & ~x[34] & ~x[37] & ~x[41] & ~x[42] & ~x[44] & ~x[46] & ~x[48] & ~x[52] & ~x[53] & ~x[54];
			partial_clause[351] 	= partial_clause_prev[351] & ~x[17];
			partial_clause[352] 	= partial_clause_prev[352] & 1'b1;
			partial_clause[353] 	= partial_clause_prev[353] & ~x[10];
			partial_clause[354] 	= partial_clause_prev[354] & ~x[13] & ~x[23];
			partial_clause[355] 	= partial_clause_prev[355] & 1'b1;
			partial_clause[356] 	= partial_clause_prev[356] & ~x[29] & ~x[41];
			partial_clause[357] 	= partial_clause_prev[357] & 1'b1;
			partial_clause[358] 	= partial_clause_prev[358] & ~x[4] & ~x[5] & ~x[7] & ~x[9] & ~x[10] & ~x[18] & ~x[21] & ~x[27] & ~x[31] & ~x[34] & ~x[38] & ~x[39] & ~x[41] & ~x[45];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[27] & ~x[39] & ~x[45];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[2] & ~x[4] & ~x[14] & ~x[16] & ~x[18] & ~x[19] & ~x[21] & ~x[27] & ~x[29] & ~x[33] & ~x[34] & ~x[39] & ~x[42] & ~x[47] & ~x[52] & ~x[54] & ~x[58] & ~x[59];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[14] & ~x[18] & ~x[22] & ~x[26] & ~x[31] & ~x[49];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[2] & ~x[8] & ~x[9] & ~x[18] & ~x[38] & ~x[39] & ~x[50];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[1] & ~x[7] & ~x[10] & ~x[16] & ~x[17] & ~x[18] & ~x[20] & ~x[28] & ~x[31] & ~x[32] & ~x[35] & ~x[41] & ~x[48] & ~x[58];
			partial_clause[364] 	= partial_clause_prev[364] & ~x[0] & ~x[27];
			partial_clause[365] 	= partial_clause_prev[365] & ~x[41];
			partial_clause[366] 	= partial_clause_prev[366] & ~x[4] & ~x[10] & ~x[11] & ~x[27] & ~x[28] & ~x[32] & ~x[33] & ~x[34] & ~x[40] & ~x[43] & ~x[44] & ~x[45] & ~x[49] & ~x[50] & ~x[54] & ~x[57] & ~x[60] & ~x[63];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[3] & ~x[5] & ~x[15] & ~x[19] & ~x[21] & ~x[24] & ~x[27] & ~x[45] & ~x[59];
			partial_clause[368] 	= partial_clause_prev[368] & 1'b1;
			partial_clause[369] 	= partial_clause_prev[369] & ~x[37] & ~x[47];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[6] & ~x[20] & ~x[34] & ~x[36] & ~x[41] & ~x[47] & ~x[58];
			partial_clause[371] 	= partial_clause_prev[371] & 1'b1;
			partial_clause[372] 	= partial_clause_prev[372] & ~x[1] & ~x[3] & ~x[9] & ~x[15] & ~x[19] & ~x[38] & ~x[44] & ~x[55] & ~x[61] & ~x[63];
			partial_clause[373] 	= partial_clause_prev[373] & ~x[28] & ~x[37];
			partial_clause[374] 	= partial_clause_prev[374] & ~x[0] & ~x[10] & ~x[34] & ~x[38] & ~x[45] & ~x[46];
			partial_clause[375] 	= partial_clause_prev[375] & ~x[37] & ~x[58];
			partial_clause[376] 	= partial_clause_prev[376] & ~x[0] & ~x[1] & ~x[5] & ~x[9] & ~x[23] & ~x[36] & ~x[37] & ~x[44] & ~x[47] & ~x[52] & ~x[54] & ~x[55];
			partial_clause[377] 	= partial_clause_prev[377] & ~x[2] & ~x[7] & ~x[8] & ~x[12] & ~x[16] & ~x[18] & ~x[25] & ~x[26] & ~x[36] & ~x[37] & ~x[39] & ~x[42] & ~x[48];
			partial_clause[378] 	= partial_clause_prev[378] & ~x[12] & ~x[46];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[3] & ~x[18] & ~x[27] & ~x[33];
			partial_clause[380] 	= partial_clause_prev[380] & 1'b1;
			partial_clause[381] 	= partial_clause_prev[381] & ~x[1] & ~x[11] & ~x[12] & ~x[14] & ~x[17] & ~x[23] & ~x[25] & ~x[26] & ~x[42] & ~x[43] & ~x[44] & ~x[47] & ~x[50] & ~x[54];
			partial_clause[382] 	= partial_clause_prev[382] & 1'b1;
			partial_clause[383] 	= partial_clause_prev[383] & ~x[36];
			partial_clause[384] 	= partial_clause_prev[384] & 1'b1;
			partial_clause[385] 	= partial_clause_prev[385] & 1'b1;
			partial_clause[386] 	= partial_clause_prev[386] & ~x[8];
			partial_clause[387] 	= partial_clause_prev[387] & ~x[0] & ~x[3] & ~x[5] & ~x[6] & ~x[9] & ~x[19] & ~x[20] & ~x[21] & ~x[24] & ~x[25] & ~x[27] & ~x[31] & ~x[34] & ~x[40] & ~x[44] & ~x[50] & ~x[53] & ~x[54] & ~x[56];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[2] & ~x[6] & ~x[9] & ~x[10] & ~x[11] & ~x[14] & ~x[19] & ~x[21] & ~x[25] & ~x[32] & ~x[33] & ~x[36] & ~x[44] & ~x[49] & ~x[54] & ~x[55] & ~x[57];
			partial_clause[389] 	= partial_clause_prev[389] & 1'b1;
			partial_clause[390] 	= partial_clause_prev[390] & ~x[2] & ~x[3] & ~x[11] & ~x[21] & ~x[25] & ~x[26] & ~x[33] & ~x[36] & ~x[39] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[50] & ~x[54];
			partial_clause[391] 	= partial_clause_prev[391] & 1'b1;
			partial_clause[392] 	= partial_clause_prev[392] & 1'b1;
			partial_clause[393] 	= partial_clause_prev[393] & 1'b1;
			partial_clause[394] 	= partial_clause_prev[394] & ~x[9] & ~x[17] & ~x[37] & ~x[39];
			partial_clause[395] 	= partial_clause_prev[395] & 1'b1;
			partial_clause[396] 	= partial_clause_prev[396] & 1'b1;
			partial_clause[397] 	= partial_clause_prev[397] & ~x[48];
			partial_clause[398] 	= partial_clause_prev[398] & 1'b1;
			partial_clause[399] 	= partial_clause_prev[399] & 1'b1;
			partial_clause[400] 	= partial_clause_prev[400] & ~x[2] & ~x[3] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[19] & ~x[25] & ~x[29] & ~x[32] & ~x[55] & ~x[57] & ~x[58] & ~x[59];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[1] & ~x[7] & ~x[10] & ~x[16] & ~x[31] & ~x[40] & ~x[42] & ~x[50] & ~x[53];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[1] & ~x[3] & ~x[4] & ~x[6] & ~x[10] & ~x[16] & ~x[18] & ~x[46] & ~x[48] & ~x[56] & ~x[61];
			partial_clause[403] 	= partial_clause_prev[403] & ~x[45];
			partial_clause[404] 	= partial_clause_prev[404] & 1'b1;
			partial_clause[405] 	= partial_clause_prev[405] & ~x[3] & ~x[8] & ~x[10] & ~x[35] & ~x[38] & ~x[43] & ~x[62];
			partial_clause[406] 	= partial_clause_prev[406] & ~x[2] & ~x[9] & ~x[20] & ~x[22] & ~x[23] & ~x[25] & ~x[35] & ~x[44] & ~x[52];
			partial_clause[407] 	= partial_clause_prev[407] & ~x[14] & ~x[23];
			partial_clause[408] 	= partial_clause_prev[408] & ~x[15] & ~x[35] & ~x[58] & ~x[63];
			partial_clause[409] 	= partial_clause_prev[409] & ~x[3] & ~x[7] & ~x[8] & ~x[9] & ~x[11] & ~x[14] & ~x[18] & ~x[19] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & ~x[28] & ~x[30] & ~x[34] & ~x[38] & ~x[41] & ~x[43] & ~x[44] & ~x[46] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[53] & ~x[54] & ~x[55] & ~x[57];
			partial_clause[410] 	= partial_clause_prev[410] & ~x[14] & ~x[18] & ~x[29] & ~x[42] & ~x[43] & ~x[51] & ~x[61];
			partial_clause[411] 	= partial_clause_prev[411] & ~x[6] & ~x[8] & ~x[22] & ~x[35] & ~x[40] & ~x[50];
			partial_clause[412] 	= partial_clause_prev[412] & ~x[0] & ~x[6] & ~x[9] & ~x[10] & ~x[15] & ~x[18] & ~x[21] & ~x[43] & ~x[46] & ~x[48] & ~x[50] & ~x[57] & ~x[62];
			partial_clause[413] 	= partial_clause_prev[413] & ~x[11] & ~x[33] & ~x[43] & ~x[54] & ~x[57];
			partial_clause[414] 	= partial_clause_prev[414] & ~x[0] & ~x[15] & ~x[17] & ~x[24] & ~x[27] & ~x[32] & ~x[33] & ~x[38] & ~x[39] & ~x[44] & ~x[51] & ~x[58] & ~x[60];
			partial_clause[415] 	= partial_clause_prev[415] & ~x[6] & ~x[32] & ~x[50];
			partial_clause[416] 	= partial_clause_prev[416] & ~x[0] & ~x[9] & ~x[13] & ~x[22] & ~x[45] & ~x[46] & ~x[47] & ~x[51] & ~x[53] & ~x[55] & ~x[57] & ~x[60];
			partial_clause[417] 	= partial_clause_prev[417] & ~x[23] & ~x[29];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[0] & ~x[1] & ~x[4] & ~x[13] & ~x[15] & ~x[21] & ~x[22] & ~x[24] & ~x[25] & ~x[29] & ~x[45] & ~x[48] & ~x[53] & ~x[54] & ~x[56];
			partial_clause[419] 	= partial_clause_prev[419] & 1'b1;
			partial_clause[420] 	= partial_clause_prev[420] & ~x[42] & ~x[49];
			partial_clause[421] 	= partial_clause_prev[421] & ~x[8] & ~x[10] & ~x[14] & ~x[18] & ~x[24] & ~x[27] & ~x[32] & ~x[34] & ~x[37] & ~x[41] & ~x[43] & ~x[51] & ~x[57] & ~x[60] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[422] 	= partial_clause_prev[422] & ~x[1] & ~x[2] & ~x[12] & ~x[19] & ~x[31] & ~x[35] & ~x[36] & ~x[41] & ~x[61];
			partial_clause[423] 	= partial_clause_prev[423] & ~x[1] & ~x[7] & ~x[40] & ~x[42] & ~x[47] & ~x[52];
			partial_clause[424] 	= partial_clause_prev[424] & ~x[10] & ~x[51] & ~x[60];
			partial_clause[425] 	= partial_clause_prev[425] & 1'b1;
			partial_clause[426] 	= partial_clause_prev[426] & ~x[0] & ~x[1] & ~x[5] & ~x[7] & ~x[8] & ~x[11] & ~x[14] & ~x[15] & ~x[16] & ~x[23] & ~x[26] & ~x[34] & ~x[35] & ~x[39] & ~x[40] & ~x[41] & ~x[52] & ~x[53] & ~x[54] & ~x[58] & ~x[60] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[0] & ~x[12] & ~x[21] & ~x[34] & ~x[43] & ~x[47] & ~x[50] & ~x[54] & ~x[56] & ~x[61];
			partial_clause[428] 	= partial_clause_prev[428] & ~x[16];
			partial_clause[429] 	= partial_clause_prev[429] & 1'b1;
			partial_clause[430] 	= partial_clause_prev[430] & ~x[6] & ~x[10] & ~x[16] & ~x[22] & ~x[23] & ~x[31] & ~x[37] & ~x[46] & ~x[52] & ~x[53];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[8];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[6] & ~x[9] & ~x[11] & ~x[12] & ~x[14] & ~x[17] & ~x[21] & ~x[23] & ~x[30] & ~x[43] & ~x[44] & ~x[46] & ~x[51] & ~x[55] & ~x[57];
			partial_clause[433] 	= partial_clause_prev[433] & ~x[42];
			partial_clause[434] 	= partial_clause_prev[434] & ~x[33];
			partial_clause[435] 	= partial_clause_prev[435] & ~x[0] & ~x[7] & ~x[11] & ~x[12] & ~x[15] & ~x[19] & ~x[25] & ~x[27] & ~x[28] & ~x[31] & ~x[32] & ~x[33] & ~x[36] & ~x[37] & ~x[43] & ~x[44] & ~x[47] & ~x[50] & ~x[51] & ~x[53] & ~x[55] & ~x[56] & ~x[57];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[8] & ~x[25] & ~x[39] & ~x[44] & ~x[51];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[7] & ~x[9] & ~x[12] & ~x[13] & ~x[23] & ~x[25] & ~x[37] & ~x[39] & ~x[40] & ~x[43] & ~x[44] & ~x[45] & ~x[46] & ~x[50] & ~x[52] & ~x[53] & ~x[54] & ~x[63];
			partial_clause[438] 	= partial_clause_prev[438] & ~x[24] & ~x[52];
			partial_clause[439] 	= partial_clause_prev[439] & ~x[15] & ~x[16] & ~x[19] & ~x[21] & ~x[24] & ~x[25] & ~x[48];
			partial_clause[440] 	= partial_clause_prev[440] & 1'b1;
			partial_clause[441] 	= partial_clause_prev[441] & ~x[2] & ~x[18] & ~x[33] & ~x[35] & ~x[46];
			partial_clause[442] 	= partial_clause_prev[442] & 1'b1;
			partial_clause[443] 	= partial_clause_prev[443] & ~x[0] & ~x[3] & ~x[6] & ~x[8] & ~x[11] & ~x[24] & ~x[35] & ~x[36] & ~x[38] & ~x[39] & ~x[41] & ~x[46] & ~x[53];
			partial_clause[444] 	= partial_clause_prev[444] & 1'b1;
			partial_clause[445] 	= partial_clause_prev[445] & ~x[62];
			partial_clause[446] 	= partial_clause_prev[446] & ~x[16] & ~x[19] & ~x[25] & ~x[28] & ~x[29] & ~x[33] & ~x[37] & ~x[42] & ~x[43] & ~x[45] & ~x[46] & ~x[54];
			partial_clause[447] 	= partial_clause_prev[447] & ~x[10] & ~x[11] & ~x[13] & ~x[22] & ~x[25] & ~x[27] & ~x[36] & ~x[37] & ~x[38];
			partial_clause[448] 	= partial_clause_prev[448] & 1'b1;
			partial_clause[449] 	= partial_clause_prev[449] & ~x[1] & ~x[20] & ~x[27] & ~x[29] & ~x[45] & ~x[52] & ~x[54];
			partial_clause[450] 	= partial_clause_prev[450] & ~x[26] & ~x[33] & ~x[49] & ~x[56];
			partial_clause[451] 	= partial_clause_prev[451] & 1'b1;
			partial_clause[452] 	= partial_clause_prev[452] & 1'b1;
			partial_clause[453] 	= partial_clause_prev[453] & ~x[42] & ~x[44];
			partial_clause[454] 	= partial_clause_prev[454] & ~x[34] & ~x[57];
			partial_clause[455] 	= partial_clause_prev[455] & ~x[0] & ~x[20] & ~x[21] & ~x[23] & ~x[28] & ~x[36] & ~x[53] & ~x[55] & ~x[59];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[14] & ~x[18] & ~x[22] & ~x[24] & ~x[26] & ~x[30] & ~x[32] & ~x[40] & ~x[41] & ~x[44] & ~x[46] & ~x[50] & ~x[57] & ~x[58];
			partial_clause[457] 	= partial_clause_prev[457] & 1'b1;
			partial_clause[458] 	= partial_clause_prev[458] & ~x[0] & ~x[10] & ~x[13] & ~x[16] & ~x[17] & ~x[29] & ~x[41] & ~x[45] & ~x[47] & ~x[54];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[5] & ~x[6] & ~x[9] & ~x[10] & ~x[21] & ~x[43];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[5] & ~x[7] & ~x[12] & ~x[19] & ~x[24] & ~x[31] & ~x[34] & ~x[36] & ~x[41] & ~x[44] & ~x[45] & ~x[60];
			partial_clause[461] 	= partial_clause_prev[461] & ~x[0] & ~x[2] & ~x[15] & ~x[21] & ~x[23] & ~x[24] & ~x[28] & ~x[35] & ~x[38] & ~x[61];
			partial_clause[462] 	= partial_clause_prev[462] & ~x[12] & ~x[22] & ~x[25];
			partial_clause[463] 	= partial_clause_prev[463] & ~x[57];
			partial_clause[464] 	= partial_clause_prev[464] & ~x[10] & ~x[13] & ~x[15] & ~x[16] & ~x[20] & ~x[26] & ~x[28] & ~x[33] & ~x[35] & ~x[38] & ~x[40] & ~x[57];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[6] & ~x[8] & ~x[14] & ~x[25] & ~x[27] & ~x[40] & ~x[48] & ~x[52] & ~x[55];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[10] & ~x[11] & ~x[16] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[23] & ~x[27] & ~x[34] & ~x[39] & ~x[40] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[55] & ~x[56];
			partial_clause[467] 	= partial_clause_prev[467] & ~x[24] & ~x[25] & ~x[31] & ~x[52];
			partial_clause[468] 	= partial_clause_prev[468] & ~x[4] & ~x[12] & ~x[14] & ~x[16] & ~x[19];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[9] & ~x[11] & ~x[13] & ~x[18] & ~x[24] & ~x[28] & ~x[36] & ~x[49] & ~x[55];
			partial_clause[470] 	= partial_clause_prev[470] & ~x[38] & ~x[45];
			partial_clause[471] 	= partial_clause_prev[471] & ~x[1] & ~x[3] & ~x[6] & ~x[22] & ~x[28] & ~x[32] & ~x[44] & ~x[50] & ~x[54];
			partial_clause[472] 	= partial_clause_prev[472] & ~x[21] & ~x[35] & ~x[59];
			partial_clause[473] 	= partial_clause_prev[473] & ~x[6] & ~x[10] & ~x[14] & ~x[18] & ~x[28] & ~x[29] & ~x[30] & ~x[35] & ~x[36] & ~x[37] & ~x[42] & ~x[44] & ~x[46] & ~x[54];
			partial_clause[474] 	= partial_clause_prev[474] & 1'b1;
			partial_clause[475] 	= partial_clause_prev[475] & ~x[16] & ~x[20] & ~x[26] & ~x[34] & ~x[42] & ~x[44] & ~x[62];
			partial_clause[476] 	= partial_clause_prev[476] & ~x[48];
			partial_clause[477] 	= partial_clause_prev[477] & ~x[18] & ~x[24] & ~x[43] & ~x[44];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[6] & ~x[11] & ~x[13] & ~x[16] & ~x[30] & ~x[40] & ~x[44] & ~x[47] & ~x[52];
			partial_clause[479] 	= partial_clause_prev[479] & 1'b1;
			partial_clause[480] 	= partial_clause_prev[480] & ~x[0] & ~x[1] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & ~x[30] & ~x[31] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[38] & ~x[39] & ~x[40] & ~x[42] & ~x[43] & ~x[44] & ~x[45] & ~x[46] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[54] & ~x[57];
			partial_clause[481] 	= partial_clause_prev[481] & ~x[5] & ~x[45];
			partial_clause[482] 	= partial_clause_prev[482] & ~x[5] & ~x[7] & ~x[15] & ~x[30] & ~x[49];
			partial_clause[483] 	= partial_clause_prev[483] & ~x[22];
			partial_clause[484] 	= partial_clause_prev[484] & ~x[8] & ~x[20] & ~x[47] & ~x[51];
			partial_clause[485] 	= partial_clause_prev[485] & 1'b1;
			partial_clause[486] 	= partial_clause_prev[486] & ~x[1] & ~x[3] & ~x[5] & ~x[18] & ~x[22] & ~x[23] & ~x[24] & ~x[45] & ~x[49] & ~x[52] & ~x[53] & ~x[55];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[1] & ~x[29] & ~x[49];
			partial_clause[488] 	= partial_clause_prev[488] & ~x[42];
			partial_clause[489] 	= partial_clause_prev[489] & ~x[52];
			partial_clause[490] 	= partial_clause_prev[490] & 1'b1;
			partial_clause[491] 	= partial_clause_prev[491] & 1'b1;
			partial_clause[492] 	= partial_clause_prev[492] & ~x[9] & ~x[15] & ~x[16] & ~x[26] & ~x[30] & ~x[56] & ~x[60];
			partial_clause[493] 	= partial_clause_prev[493] & ~x[30];
			partial_clause[494] 	= partial_clause_prev[494] & ~x[27] & ~x[38];
			partial_clause[495] 	= partial_clause_prev[495] & ~x[2] & ~x[4] & ~x[6] & ~x[8] & ~x[13] & ~x[15] & ~x[20] & ~x[40] & ~x[53];
			partial_clause[496] 	= partial_clause_prev[496] & 1'b1;
			partial_clause[497] 	= partial_clause_prev[497] & ~x[63];
			partial_clause[498] 	= partial_clause_prev[498] & 1'b1;
			partial_clause[499] 	= partial_clause_prev[499] & ~x[42];
		end
	end
endmodule


module HCB_2 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[3] & ~x[7] & ~x[8] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[36] & ~x[40] & ~x[41] & ~x[43];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[14] & ~x[19] & ~x[43] & ~x[48];
			partial_clause[2] 	= partial_clause_prev[2] & ~x[6];
			partial_clause[3] 	= partial_clause_prev[3] & ~x[19] & ~x[24] & ~x[41] & ~x[42];
			partial_clause[4] 	= partial_clause_prev[4] & ~x[36] & ~x[49];
			partial_clause[5] 	= partial_clause_prev[5] & ~x[10] & ~x[18] & ~x[21] & ~x[36];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[5] & x[27] & ~x[35] & ~x[37] & ~x[38] & ~x[63];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[11] & ~x[19] & ~x[38] & ~x[60];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[4] & ~x[5] & ~x[7] & ~x[9] & ~x[10] & ~x[12] & ~x[13] & ~x[14] & ~x[21] & ~x[24] & ~x[38] & ~x[44] & ~x[45];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[20] & ~x[37] & ~x[41] & ~x[62];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[1] & ~x[18] & ~x[21] & ~x[42] & ~x[43] & ~x[47] & ~x[49];
			partial_clause[11] 	= partial_clause_prev[11] & ~x[14] & ~x[39];
			partial_clause[12] 	= partial_clause_prev[12] & ~x[6] & ~x[7] & ~x[17] & ~x[33] & ~x[44];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[4] & ~x[12] & ~x[15] & ~x[16] & ~x[20] & ~x[21] & ~x[37] & ~x[39] & ~x[45];
			partial_clause[14] 	= partial_clause_prev[14] & ~x[33] & ~x[62];
			partial_clause[15] 	= partial_clause_prev[15] & 1'b1;
			partial_clause[16] 	= partial_clause_prev[16] & ~x[18] & ~x[19] & ~x[30] & ~x[46] & ~x[63];
			partial_clause[17] 	= partial_clause_prev[17] & x[54];
			partial_clause[18] 	= partial_clause_prev[18] & ~x[20] & ~x[45];
			partial_clause[19] 	= partial_clause_prev[19] & 1'b1;
			partial_clause[20] 	= partial_clause_prev[20] & ~x[8] & ~x[40];
			partial_clause[21] 	= partial_clause_prev[21] & ~x[22] & ~x[53];
			partial_clause[22] 	= partial_clause_prev[22] & ~x[49];
			partial_clause[23] 	= partial_clause_prev[23] & ~x[3] & ~x[9] & ~x[10] & ~x[12] & ~x[14] & ~x[15] & ~x[16] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[39] & ~x[40] & ~x[44];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[7] & ~x[8] & ~x[9] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[18] & ~x[34] & ~x[36] & ~x[37] & ~x[38] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[45] & ~x[46] & ~x[63];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[10] & ~x[14] & ~x[16] & ~x[20] & ~x[21] & ~x[35] & ~x[36] & ~x[37] & ~x[38] & ~x[41] & ~x[42] & ~x[43] & ~x[46] & ~x[48] & x[57];
			partial_clause[26] 	= partial_clause_prev[26] & 1'b1;
			partial_clause[27] 	= partial_clause_prev[27] & ~x[6] & ~x[12] & ~x[16] & ~x[19] & ~x[44] & ~x[46] & ~x[47] & ~x[58] & ~x[60];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[9] & ~x[20] & ~x[24] & ~x[37] & ~x[52];
			partial_clause[29] 	= partial_clause_prev[29] & ~x[1] & ~x[7] & ~x[18];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[8] & ~x[12];
			partial_clause[31] 	= partial_clause_prev[31] & ~x[16] & ~x[38] & ~x[42] & x[55];
			partial_clause[32] 	= partial_clause_prev[32] & ~x[20];
			partial_clause[33] 	= partial_clause_prev[33] & ~x[3];
			partial_clause[34] 	= partial_clause_prev[34] & ~x[3] & ~x[5] & ~x[10] & ~x[14] & ~x[16] & ~x[18] & ~x[34] & ~x[43] & ~x[45] & ~x[62];
			partial_clause[35] 	= partial_clause_prev[35] & ~x[7] & ~x[39];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[5] & ~x[38] & ~x[42] & ~x[63];
			partial_clause[37] 	= partial_clause_prev[37] & ~x[5] & ~x[14] & ~x[43] & ~x[61];
			partial_clause[38] 	= partial_clause_prev[38] & ~x[12] & ~x[13] & ~x[14] & ~x[18] & ~x[19] & ~x[44] & ~x[48];
			partial_clause[39] 	= partial_clause_prev[39] & ~x[48];
			partial_clause[40] 	= partial_clause_prev[40] & ~x[11] & ~x[40] & ~x[63];
			partial_clause[41] 	= partial_clause_prev[41] & 1'b1;
			partial_clause[42] 	= partial_clause_prev[42] & ~x[12];
			partial_clause[43] 	= partial_clause_prev[43] & ~x[18] & ~x[38] & ~x[63];
			partial_clause[44] 	= partial_clause_prev[44] & 1'b1;
			partial_clause[45] 	= partial_clause_prev[45] & ~x[63];
			partial_clause[46] 	= partial_clause_prev[46] & ~x[8] & ~x[9] & ~x[12] & ~x[17] & ~x[19] & ~x[31] & ~x[34] & ~x[36] & ~x[39] & ~x[42] & ~x[62] & ~x[63];
			partial_clause[47] 	= partial_clause_prev[47] & ~x[31] & ~x[32] & ~x[36];
			partial_clause[48] 	= partial_clause_prev[48] & 1'b1;
			partial_clause[49] 	= partial_clause_prev[49] & ~x[4];
			partial_clause[50] 	= partial_clause_prev[50] & ~x[35] & ~x[42] & ~x[44];
			partial_clause[51] 	= partial_clause_prev[51] & 1'b1;
			partial_clause[52] 	= partial_clause_prev[52] & ~x[36];
			partial_clause[53] 	= partial_clause_prev[53] & 1'b1;
			partial_clause[54] 	= partial_clause_prev[54] & 1'b1;
			partial_clause[55] 	= partial_clause_prev[55] & 1'b1;
			partial_clause[56] 	= partial_clause_prev[56] & ~x[55];
			partial_clause[57] 	= partial_clause_prev[57] & ~x[5] & ~x[18] & ~x[33];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[6] & ~x[13] & ~x[15] & ~x[40];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[2] & ~x[6] & ~x[18] & ~x[32] & ~x[34] & ~x[35] & ~x[44] & ~x[62];
			partial_clause[60] 	= partial_clause_prev[60] & 1'b1;
			partial_clause[61] 	= partial_clause_prev[61] & 1'b1;
			partial_clause[62] 	= partial_clause_prev[62] & ~x[6] & ~x[9] & ~x[12];
			partial_clause[63] 	= partial_clause_prev[63] & ~x[42];
			partial_clause[64] 	= partial_clause_prev[64] & 1'b1;
			partial_clause[65] 	= partial_clause_prev[65] & 1'b1;
			partial_clause[66] 	= partial_clause_prev[66] & 1'b1;
			partial_clause[67] 	= partial_clause_prev[67] & 1'b1;
			partial_clause[68] 	= partial_clause_prev[68] & ~x[9] & ~x[12] & ~x[37];
			partial_clause[69] 	= partial_clause_prev[69] & ~x[1] & ~x[3] & ~x[13] & ~x[14] & ~x[15] & ~x[31] & ~x[35] & ~x[38] & ~x[40] & ~x[43] & ~x[61];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[38] & ~x[46] & ~x[48];
			partial_clause[71] 	= partial_clause_prev[71] & 1'b1;
			partial_clause[72] 	= partial_clause_prev[72] & ~x[12];
			partial_clause[73] 	= partial_clause_prev[73] & 1'b1;
			partial_clause[74] 	= partial_clause_prev[74] & ~x[11] & ~x[12] & ~x[18] & ~x[38] & ~x[42] & ~x[46];
			partial_clause[75] 	= partial_clause_prev[75] & 1'b1;
			partial_clause[76] 	= partial_clause_prev[76] & ~x[6] & ~x[37] & ~x[39] & ~x[40];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[34];
			partial_clause[78] 	= partial_clause_prev[78] & ~x[12];
			partial_clause[79] 	= partial_clause_prev[79] & ~x[44] & ~x[63];
			partial_clause[80] 	= partial_clause_prev[80] & ~x[57];
			partial_clause[81] 	= partial_clause_prev[81] & 1'b1;
			partial_clause[82] 	= partial_clause_prev[82] & 1'b1;
			partial_clause[83] 	= partial_clause_prev[83] & 1'b1;
			partial_clause[84] 	= partial_clause_prev[84] & ~x[9];
			partial_clause[85] 	= partial_clause_prev[85] & ~x[4] & ~x[8] & ~x[9] & ~x[15] & ~x[34] & ~x[36] & ~x[43] & ~x[46];
			partial_clause[86] 	= partial_clause_prev[86] & 1'b1;
			partial_clause[87] 	= partial_clause_prev[87] & ~x[13] & ~x[38] & ~x[40];
			partial_clause[88] 	= partial_clause_prev[88] & ~x[16] & ~x[18] & ~x[42] & ~x[45];
			partial_clause[89] 	= partial_clause_prev[89] & 1'b1;
			partial_clause[90] 	= partial_clause_prev[90] & ~x[27];
			partial_clause[91] 	= partial_clause_prev[91] & ~x[18];
			partial_clause[92] 	= partial_clause_prev[92] & ~x[15] & ~x[20] & ~x[24] & ~x[40] & ~x[41] & ~x[52];
			partial_clause[93] 	= partial_clause_prev[93] & ~x[6] & ~x[9] & ~x[10] & ~x[16] & ~x[18] & ~x[38] & ~x[41] & ~x[46] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[94] 	= partial_clause_prev[94] & ~x[24];
			partial_clause[95] 	= partial_clause_prev[95] & ~x[9] & ~x[10] & ~x[13] & ~x[18] & ~x[20] & ~x[43] & ~x[46] & ~x[63];
			partial_clause[96] 	= partial_clause_prev[96] & ~x[27] & ~x[30];
			partial_clause[97] 	= partial_clause_prev[97] & ~x[7] & ~x[12] & ~x[14] & ~x[15] & ~x[21] & ~x[43] & ~x[48] & ~x[50];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[7] & ~x[8] & ~x[12] & ~x[19] & ~x[37] & ~x[42] & ~x[47];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[30] & ~x[31] & ~x[35] & ~x[36] & ~x[45] & ~x[46] & ~x[47];
			partial_clause[100] 	= partial_clause_prev[100] & 1'b1;
			partial_clause[101] 	= partial_clause_prev[101] & 1'b1;
			partial_clause[102] 	= partial_clause_prev[102] & ~x[0] & ~x[49];
			partial_clause[103] 	= partial_clause_prev[103] & ~x[13] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[39] & ~x[41] & ~x[43] & ~x[44] & ~x[47] & ~x[62];
			partial_clause[104] 	= partial_clause_prev[104] & ~x[3] & ~x[4] & ~x[11] & ~x[18] & ~x[61];
			partial_clause[105] 	= partial_clause_prev[105] & ~x[0] & ~x[1] & ~x[5] & ~x[10] & ~x[11] & ~x[12] & ~x[18] & ~x[34] & ~x[38] & ~x[41] & ~x[45];
			partial_clause[106] 	= partial_clause_prev[106] & ~x[13] & ~x[18] & ~x[20] & x[28] & ~x[46];
			partial_clause[107] 	= partial_clause_prev[107] & ~x[5] & ~x[11] & ~x[16] & ~x[23] & ~x[25] & ~x[32] & ~x[40] & ~x[41] & ~x[45] & ~x[63];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[5] & ~x[8] & ~x[12] & ~x[13] & ~x[17] & ~x[19] & ~x[36] & ~x[43] & ~x[46] & ~x[47] & ~x[62];
			partial_clause[109] 	= partial_clause_prev[109] & ~x[0] & ~x[54];
			partial_clause[110] 	= partial_clause_prev[110] & ~x[34];
			partial_clause[111] 	= partial_clause_prev[111] & 1'b1;
			partial_clause[112] 	= partial_clause_prev[112] & ~x[9];
			partial_clause[113] 	= partial_clause_prev[113] & ~x[26];
			partial_clause[114] 	= partial_clause_prev[114] & 1'b1;
			partial_clause[115] 	= partial_clause_prev[115] & ~x[5] & ~x[6] & ~x[15] & ~x[16] & ~x[17] & ~x[33] & ~x[38] & ~x[41] & ~x[44];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[10] & ~x[12] & ~x[43] & ~x[46] & ~x[49] & x[55] & x[56];
			partial_clause[117] 	= partial_clause_prev[117] & 1'b1;
			partial_clause[118] 	= partial_clause_prev[118] & ~x[9] & ~x[19] & ~x[39] & ~x[44] & ~x[62];
			partial_clause[119] 	= partial_clause_prev[119] & ~x[3] & ~x[6] & ~x[8] & ~x[13] & ~x[17] & ~x[32] & ~x[38] & ~x[42];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[6] & ~x[8] & ~x[9] & ~x[10] & ~x[12] & ~x[14] & ~x[18] & ~x[36] & ~x[39] & ~x[40] & ~x[44];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[9] & ~x[10] & ~x[12] & ~x[39] & ~x[41] & ~x[42] & ~x[43] & x[54];
			partial_clause[122] 	= partial_clause_prev[122] & ~x[23] & ~x[39] & ~x[50];
			partial_clause[123] 	= partial_clause_prev[123] & ~x[8] & ~x[9] & ~x[10] & ~x[13] & ~x[16] & ~x[18] & ~x[38] & ~x[40] & ~x[41] & ~x[43] & ~x[49];
			partial_clause[124] 	= partial_clause_prev[124] & 1'b1;
			partial_clause[125] 	= partial_clause_prev[125] & 1'b1;
			partial_clause[126] 	= partial_clause_prev[126] & ~x[8] & ~x[31] & ~x[34] & ~x[36] & ~x[41];
			partial_clause[127] 	= partial_clause_prev[127] & ~x[10] & ~x[12] & ~x[14] & ~x[16] & ~x[23] & ~x[35] & ~x[36] & ~x[37] & ~x[39] & ~x[44] & ~x[63];
			partial_clause[128] 	= partial_clause_prev[128] & ~x[1] & ~x[2] & ~x[22] & ~x[46];
			partial_clause[129] 	= partial_clause_prev[129] & ~x[0] & ~x[2] & ~x[10] & ~x[20] & ~x[22] & ~x[34] & ~x[42] & ~x[45] & ~x[50] & ~x[62];
			partial_clause[130] 	= partial_clause_prev[130] & ~x[4] & ~x[5] & ~x[32] & ~x[42];
			partial_clause[131] 	= partial_clause_prev[131] & ~x[14] & ~x[26] & ~x[28];
			partial_clause[132] 	= partial_clause_prev[132] & ~x[12] & ~x[14] & ~x[31] & ~x[46];
			partial_clause[133] 	= partial_clause_prev[133] & ~x[16] & ~x[20] & ~x[24];
			partial_clause[134] 	= partial_clause_prev[134] & ~x[6] & ~x[7] & ~x[20] & ~x[36] & ~x[38] & ~x[39] & ~x[41] & ~x[43] & ~x[47];
			partial_clause[135] 	= partial_clause_prev[135] & ~x[10] & ~x[41] & ~x[46];
			partial_clause[136] 	= partial_clause_prev[136] & ~x[3] & ~x[7] & ~x[8] & ~x[9] & ~x[11] & ~x[16] & ~x[42] & ~x[43] & ~x[63];
			partial_clause[137] 	= partial_clause_prev[137] & ~x[28];
			partial_clause[138] 	= partial_clause_prev[138] & ~x[13];
			partial_clause[139] 	= partial_clause_prev[139] & ~x[2] & ~x[5] & ~x[8] & ~x[10] & ~x[12] & ~x[15] & ~x[31] & ~x[43] & ~x[59];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[8] & ~x[10] & ~x[11] & ~x[13] & ~x[14] & ~x[20] & ~x[35] & ~x[38] & ~x[52] & ~x[53] & ~x[63];
			partial_clause[141] 	= partial_clause_prev[141] & ~x[20] & ~x[37] & ~x[38] & ~x[61];
			partial_clause[142] 	= partial_clause_prev[142] & ~x[5] & ~x[12] & ~x[13] & ~x[18];
			partial_clause[143] 	= partial_clause_prev[143] & ~x[41] & ~x[44] & ~x[46];
			partial_clause[144] 	= partial_clause_prev[144] & ~x[2] & ~x[10] & ~x[12] & ~x[26] & ~x[27] & ~x[28] & ~x[30] & ~x[39] & ~x[41] & ~x[42] & ~x[43] & ~x[47];
			partial_clause[145] 	= partial_clause_prev[145] & ~x[45];
			partial_clause[146] 	= partial_clause_prev[146] & ~x[13] & ~x[44];
			partial_clause[147] 	= partial_clause_prev[147] & ~x[13] & ~x[47];
			partial_clause[148] 	= partial_clause_prev[148] & ~x[4] & ~x[15] & ~x[18] & ~x[36];
			partial_clause[149] 	= partial_clause_prev[149] & ~x[17] & ~x[29] & ~x[56] & ~x[57];
			partial_clause[150] 	= partial_clause_prev[150] & ~x[13] & ~x[15];
			partial_clause[151] 	= partial_clause_prev[151] & 1'b1;
			partial_clause[152] 	= partial_clause_prev[152] & ~x[15];
			partial_clause[153] 	= partial_clause_prev[153] & ~x[11] & ~x[12] & ~x[39] & ~x[41] & ~x[62];
			partial_clause[154] 	= partial_clause_prev[154] & 1'b1;
			partial_clause[155] 	= partial_clause_prev[155] & 1'b1;
			partial_clause[156] 	= partial_clause_prev[156] & ~x[10];
			partial_clause[157] 	= partial_clause_prev[157] & 1'b1;
			partial_clause[158] 	= partial_clause_prev[158] & ~x[9] & ~x[11] & ~x[12] & ~x[14] & ~x[16] & ~x[19] & ~x[20] & ~x[22] & ~x[24] & ~x[37] & ~x[38] & ~x[45] & ~x[46];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[8] & ~x[9] & ~x[10] & ~x[17] & ~x[44];
			partial_clause[160] 	= partial_clause_prev[160] & ~x[6];
			partial_clause[161] 	= partial_clause_prev[161] & ~x[8] & ~x[15] & ~x[30] & ~x[38] & ~x[45];
			partial_clause[162] 	= partial_clause_prev[162] & ~x[7] & ~x[15] & ~x[16] & ~x[20] & ~x[35] & ~x[38];
			partial_clause[163] 	= partial_clause_prev[163] & 1'b1;
			partial_clause[164] 	= partial_clause_prev[164] & ~x[22] & ~x[43];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[2] & ~x[15] & ~x[20] & ~x[22] & ~x[25] & ~x[32] & ~x[35] & ~x[38] & ~x[43];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[5] & ~x[7] & ~x[9] & ~x[15] & ~x[45] & ~x[63];
			partial_clause[167] 	= partial_clause_prev[167] & x[28];
			partial_clause[168] 	= partial_clause_prev[168] & ~x[10];
			partial_clause[169] 	= partial_clause_prev[169] & 1'b1;
			partial_clause[170] 	= partial_clause_prev[170] & ~x[24] & ~x[52];
			partial_clause[171] 	= partial_clause_prev[171] & ~x[0] & ~x[11];
			partial_clause[172] 	= partial_clause_prev[172] & ~x[26] & ~x[53];
			partial_clause[173] 	= partial_clause_prev[173] & ~x[11] & ~x[13] & ~x[21] & ~x[36] & ~x[38] & ~x[42] & x[58];
			partial_clause[174] 	= partial_clause_prev[174] & ~x[3] & ~x[30];
			partial_clause[175] 	= partial_clause_prev[175] & ~x[56];
			partial_clause[176] 	= partial_clause_prev[176] & ~x[17];
			partial_clause[177] 	= partial_clause_prev[177] & ~x[15] & ~x[26] & ~x[27] & ~x[36] & ~x[38] & ~x[40] & ~x[63];
			partial_clause[178] 	= partial_clause_prev[178] & ~x[3] & ~x[17] & ~x[42];
			partial_clause[179] 	= partial_clause_prev[179] & ~x[55];
			partial_clause[180] 	= partial_clause_prev[180] & ~x[10];
			partial_clause[181] 	= partial_clause_prev[181] & 1'b1;
			partial_clause[182] 	= partial_clause_prev[182] & ~x[27];
			partial_clause[183] 	= partial_clause_prev[183] & ~x[3] & ~x[13] & ~x[14] & ~x[16] & ~x[23] & ~x[37] & ~x[44] & ~x[45] & ~x[50];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[12] & ~x[15] & ~x[16] & ~x[17] & ~x[20] & ~x[25] & ~x[38] & ~x[39] & ~x[41] & ~x[46];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[10] & ~x[63];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[9] & ~x[20] & ~x[22] & ~x[35] & ~x[39] & ~x[42] & ~x[43] & ~x[46] & ~x[62];
			partial_clause[187] 	= partial_clause_prev[187] & ~x[7] & ~x[8] & ~x[12] & ~x[34] & ~x[35] & ~x[42] & ~x[59] & ~x[61];
			partial_clause[188] 	= partial_clause_prev[188] & ~x[34];
			partial_clause[189] 	= partial_clause_prev[189] & 1'b1;
			partial_clause[190] 	= partial_clause_prev[190] & ~x[7] & ~x[17] & ~x[19] & ~x[24] & ~x[26] & ~x[46];
			partial_clause[191] 	= partial_clause_prev[191] & 1'b1;
			partial_clause[192] 	= partial_clause_prev[192] & ~x[11] & ~x[13] & ~x[34];
			partial_clause[193] 	= partial_clause_prev[193] & ~x[8] & ~x[9] & ~x[29] & ~x[43] & ~x[48] & ~x[60];
			partial_clause[194] 	= partial_clause_prev[194] & ~x[11] & x[59];
			partial_clause[195] 	= partial_clause_prev[195] & ~x[7] & ~x[12] & ~x[15] & ~x[31] & ~x[33] & ~x[35] & ~x[36] & ~x[43];
			partial_clause[196] 	= partial_clause_prev[196] & ~x[6] & ~x[26] & ~x[38];
			partial_clause[197] 	= partial_clause_prev[197] & ~x[9] & ~x[11] & ~x[13] & ~x[14] & ~x[38] & ~x[49];
			partial_clause[198] 	= partial_clause_prev[198] & ~x[29];
			partial_clause[199] 	= partial_clause_prev[199] & 1'b1;
			partial_clause[200] 	= partial_clause_prev[200] & 1'b1;
			partial_clause[201] 	= partial_clause_prev[201] & ~x[7] & ~x[13] & ~x[38];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[8] & ~x[9] & ~x[13] & ~x[16] & ~x[17] & ~x[20] & ~x[33] & ~x[37] & ~x[38] & ~x[39] & ~x[49] & ~x[62];
			partial_clause[203] 	= partial_clause_prev[203] & 1'b1;
			partial_clause[204] 	= partial_clause_prev[204] & ~x[0] & ~x[10] & ~x[11] & ~x[14] & ~x[15] & ~x[21] & ~x[22] & ~x[32] & ~x[43] & ~x[50];
			partial_clause[205] 	= partial_clause_prev[205] & ~x[4] & ~x[28];
			partial_clause[206] 	= partial_clause_prev[206] & ~x[7] & ~x[13] & ~x[15] & ~x[35] & ~x[43];
			partial_clause[207] 	= partial_clause_prev[207] & ~x[11] & ~x[12] & ~x[20] & ~x[33] & ~x[41] & ~x[45] & ~x[61];
			partial_clause[208] 	= partial_clause_prev[208] & ~x[0] & ~x[6] & ~x[26];
			partial_clause[209] 	= partial_clause_prev[209] & ~x[51];
			partial_clause[210] 	= partial_clause_prev[210] & ~x[18] & ~x[39] & ~x[45];
			partial_clause[211] 	= partial_clause_prev[211] & ~x[39];
			partial_clause[212] 	= partial_clause_prev[212] & ~x[12] & ~x[21] & ~x[41] & ~x[53];
			partial_clause[213] 	= partial_clause_prev[213] & 1'b1;
			partial_clause[214] 	= partial_clause_prev[214] & ~x[7];
			partial_clause[215] 	= partial_clause_prev[215] & ~x[42];
			partial_clause[216] 	= partial_clause_prev[216] & x[59];
			partial_clause[217] 	= partial_clause_prev[217] & ~x[8] & ~x[13] & ~x[14] & ~x[46];
			partial_clause[218] 	= partial_clause_prev[218] & ~x[44];
			partial_clause[219] 	= partial_clause_prev[219] & ~x[61];
			partial_clause[220] 	= partial_clause_prev[220] & ~x[0] & ~x[1] & ~x[7] & ~x[8] & ~x[16] & ~x[17] & ~x[20] & ~x[24] & ~x[25] & ~x[28] & ~x[29] & ~x[33] & ~x[34] & ~x[36] & ~x[40] & ~x[41] & ~x[50] & ~x[53] & ~x[55];
			partial_clause[221] 	= partial_clause_prev[221] & ~x[10] & ~x[23] & ~x[25] & ~x[29] & ~x[37];
			partial_clause[222] 	= partial_clause_prev[222] & 1'b1;
			partial_clause[223] 	= partial_clause_prev[223] & ~x[1] & ~x[2] & ~x[46];
			partial_clause[224] 	= partial_clause_prev[224] & ~x[15] & ~x[20] & ~x[39] & ~x[43] & ~x[44] & ~x[46] & ~x[49];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[17] & x[28];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[14] & ~x[16] & ~x[17] & ~x[19] & ~x[22] & ~x[37] & ~x[39] & ~x[42] & ~x[45] & ~x[47] & ~x[48] & ~x[49];
			partial_clause[227] 	= partial_clause_prev[227] & 1'b1;
			partial_clause[228] 	= partial_clause_prev[228] & ~x[12] & ~x[17] & ~x[44] & ~x[47] & ~x[50];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[21] & ~x[35] & ~x[36] & ~x[41] & ~x[44] & ~x[47] & ~x[49] & ~x[63];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[1] & ~x[2] & ~x[3] & ~x[7] & ~x[9] & ~x[14] & ~x[17] & ~x[18] & ~x[33] & ~x[40] & ~x[43] & ~x[46];
			partial_clause[231] 	= partial_clause_prev[231] & ~x[9] & ~x[15] & x[29] & ~x[40];
			partial_clause[232] 	= partial_clause_prev[232] & 1'b1;
			partial_clause[233] 	= partial_clause_prev[233] & ~x[8] & ~x[10] & ~x[37] & x[54] & ~x[63];
			partial_clause[234] 	= partial_clause_prev[234] & ~x[38] & ~x[60];
			partial_clause[235] 	= partial_clause_prev[235] & 1'b1;
			partial_clause[236] 	= partial_clause_prev[236] & ~x[14];
			partial_clause[237] 	= partial_clause_prev[237] & ~x[19] & ~x[21];
			partial_clause[238] 	= partial_clause_prev[238] & ~x[21] & ~x[35] & ~x[40] & ~x[52];
			partial_clause[239] 	= partial_clause_prev[239] & ~x[35];
			partial_clause[240] 	= partial_clause_prev[240] & ~x[8] & ~x[15] & ~x[17] & ~x[20] & ~x[38] & ~x[39] & ~x[49];
			partial_clause[241] 	= partial_clause_prev[241] & ~x[37] & ~x[42];
			partial_clause[242] 	= partial_clause_prev[242] & ~x[12] & ~x[15] & ~x[42] & ~x[47] & ~x[48] & ~x[54];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[5] & ~x[38] & ~x[39] & ~x[42] & ~x[43] & ~x[62] & ~x[63];
			partial_clause[244] 	= partial_clause_prev[244] & ~x[26];
			partial_clause[245] 	= partial_clause_prev[245] & 1'b1;
			partial_clause[246] 	= partial_clause_prev[246] & ~x[41] & x[52] & ~x[62];
			partial_clause[247] 	= partial_clause_prev[247] & ~x[9] & ~x[12] & ~x[18] & ~x[39] & ~x[40] & ~x[45] & ~x[47] & ~x[48];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[10] & ~x[11] & ~x[13] & ~x[15] & ~x[16] & ~x[30] & ~x[36] & ~x[37] & ~x[39] & ~x[41] & ~x[44] & ~x[63];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[8] & ~x[33] & ~x[37];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[4] & ~x[5] & ~x[7] & ~x[9] & ~x[11] & ~x[35] & ~x[37] & ~x[39] & ~x[40] & ~x[41] & ~x[47];
			partial_clause[251] 	= partial_clause_prev[251] & ~x[5] & ~x[23];
			partial_clause[252] 	= partial_clause_prev[252] & ~x[9] & ~x[11] & ~x[13] & ~x[16] & ~x[17] & ~x[18] & ~x[33] & ~x[34] & ~x[38] & ~x[39] & ~x[40] & ~x[42] & ~x[43] & ~x[45] & ~x[46] & ~x[59];
			partial_clause[253] 	= partial_clause_prev[253] & ~x[15] & ~x[34] & ~x[35];
			partial_clause[254] 	= partial_clause_prev[254] & ~x[17] & ~x[40] & x[55];
			partial_clause[255] 	= partial_clause_prev[255] & ~x[8] & ~x[12] & ~x[13] & ~x[14] & ~x[15];
			partial_clause[256] 	= partial_clause_prev[256] & 1'b1;
			partial_clause[257] 	= partial_clause_prev[257] & ~x[3] & ~x[14] & ~x[21] & ~x[63];
			partial_clause[258] 	= partial_clause_prev[258] & ~x[1] & ~x[46];
			partial_clause[259] 	= partial_clause_prev[259] & 1'b1;
			partial_clause[260] 	= partial_clause_prev[260] & ~x[9] & ~x[10] & ~x[42] & ~x[63];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[7] & ~x[12] & ~x[17] & ~x[20] & ~x[36] & ~x[38] & ~x[39] & ~x[40] & ~x[44];
			partial_clause[262] 	= partial_clause_prev[262] & ~x[6] & ~x[35] & ~x[36] & ~x[41];
			partial_clause[263] 	= partial_clause_prev[263] & 1'b1;
			partial_clause[264] 	= partial_clause_prev[264] & ~x[17] & ~x[35] & ~x[40];
			partial_clause[265] 	= partial_clause_prev[265] & 1'b1;
			partial_clause[266] 	= partial_clause_prev[266] & ~x[0] & ~x[7] & ~x[8] & ~x[13] & ~x[34] & ~x[39] & ~x[41];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[1] & ~x[5] & ~x[7] & ~x[9] & ~x[14] & ~x[16] & ~x[17] & ~x[18] & ~x[23] & ~x[30] & ~x[34] & ~x[41] & ~x[42] & ~x[46];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[16] & ~x[18] & ~x[38];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[8] & ~x[9] & ~x[11] & ~x[12] & ~x[14] & ~x[15] & ~x[16] & ~x[19] & ~x[21] & ~x[36] & ~x[37] & ~x[38] & ~x[40] & ~x[41] & ~x[43] & ~x[44] & ~x[45] & ~x[48];
			partial_clause[270] 	= partial_clause_prev[270] & 1'b1;
			partial_clause[271] 	= partial_clause_prev[271] & 1'b1;
			partial_clause[272] 	= partial_clause_prev[272] & ~x[10] & ~x[36] & ~x[38] & ~x[44];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[5] & ~x[9] & ~x[10] & ~x[16] & ~x[18] & ~x[20] & ~x[38] & ~x[39] & ~x[43] & ~x[45];
			partial_clause[274] 	= partial_clause_prev[274] & ~x[7] & ~x[13] & ~x[15] & x[25] & ~x[39] & ~x[42];
			partial_clause[275] 	= partial_clause_prev[275] & ~x[18] & ~x[22] & ~x[40] & ~x[42];
			partial_clause[276] 	= partial_clause_prev[276] & ~x[7] & ~x[16] & ~x[23] & ~x[40];
			partial_clause[277] 	= partial_clause_prev[277] & ~x[24] & ~x[44] & ~x[48] & ~x[50];
			partial_clause[278] 	= partial_clause_prev[278] & 1'b1;
			partial_clause[279] 	= partial_clause_prev[279] & ~x[7] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[17] & ~x[20] & ~x[22] & ~x[40] & ~x[45] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[280] 	= partial_clause_prev[280] & 1'b1;
			partial_clause[281] 	= partial_clause_prev[281] & ~x[6] & ~x[8] & ~x[12] & ~x[16] & ~x[17] & ~x[20] & ~x[43] & ~x[47] & ~x[50] & ~x[63];
			partial_clause[282] 	= partial_clause_prev[282] & ~x[7] & ~x[14] & ~x[35] & ~x[39] & x[55];
			partial_clause[283] 	= partial_clause_prev[283] & 1'b1;
			partial_clause[284] 	= partial_clause_prev[284] & ~x[36];
			partial_clause[285] 	= partial_clause_prev[285] & 1'b1;
			partial_clause[286] 	= partial_clause_prev[286] & ~x[1] & ~x[24] & ~x[27] & ~x[48];
			partial_clause[287] 	= partial_clause_prev[287] & ~x[9] & ~x[12] & ~x[36] & ~x[40] & ~x[41] & ~x[43];
			partial_clause[288] 	= partial_clause_prev[288] & ~x[26] & ~x[30] & ~x[53] & ~x[60];
			partial_clause[289] 	= partial_clause_prev[289] & ~x[9] & ~x[10] & ~x[35] & x[51] & ~x[60] & ~x[61];
			partial_clause[290] 	= partial_clause_prev[290] & ~x[7] & ~x[35];
			partial_clause[291] 	= partial_clause_prev[291] & ~x[24] & ~x[52];
			partial_clause[292] 	= partial_clause_prev[292] & ~x[0] & ~x[11] & ~x[27] & ~x[38];
			partial_clause[293] 	= partial_clause_prev[293] & ~x[2] & ~x[34] & ~x[36];
			partial_clause[294] 	= partial_clause_prev[294] & ~x[3] & ~x[8] & ~x[23];
			partial_clause[295] 	= partial_clause_prev[295] & ~x[17] & ~x[19] & ~x[36];
			partial_clause[296] 	= partial_clause_prev[296] & ~x[54];
			partial_clause[297] 	= partial_clause_prev[297] & ~x[10] & ~x[11] & ~x[16] & ~x[22];
			partial_clause[298] 	= partial_clause_prev[298] & 1'b1;
			partial_clause[299] 	= partial_clause_prev[299] & ~x[5] & ~x[7] & ~x[13] & ~x[36] & ~x[38] & ~x[39] & ~x[48];
			partial_clause[300] 	= partial_clause_prev[300] & ~x[11] & ~x[12] & ~x[21] & x[27];
			partial_clause[301] 	= partial_clause_prev[301] & ~x[1] & ~x[6] & ~x[7] & ~x[12] & ~x[18] & ~x[46] & ~x[63];
			partial_clause[302] 	= partial_clause_prev[302] & ~x[40];
			partial_clause[303] 	= partial_clause_prev[303] & ~x[23] & ~x[43] & ~x[47] & ~x[48];
			partial_clause[304] 	= partial_clause_prev[304] & ~x[7] & ~x[38];
			partial_clause[305] 	= partial_clause_prev[305] & ~x[12] & ~x[15] & ~x[47];
			partial_clause[306] 	= partial_clause_prev[306] & ~x[14] & ~x[15] & ~x[16];
			partial_clause[307] 	= partial_clause_prev[307] & ~x[5] & ~x[10] & ~x[12] & ~x[21] & ~x[43] & ~x[44];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[9] & ~x[11] & ~x[29] & ~x[37] & ~x[43] & ~x[63];
			partial_clause[309] 	= partial_clause_prev[309] & ~x[17] & ~x[20] & ~x[38];
			partial_clause[310] 	= partial_clause_prev[310] & 1'b1;
			partial_clause[311] 	= partial_clause_prev[311] & ~x[27];
			partial_clause[312] 	= partial_clause_prev[312] & ~x[45] & ~x[47];
			partial_clause[313] 	= partial_clause_prev[313] & 1'b1;
			partial_clause[314] 	= partial_clause_prev[314] & ~x[3];
			partial_clause[315] 	= partial_clause_prev[315] & ~x[2] & ~x[24] & ~x[29] & ~x[46] & ~x[48] & ~x[50] & ~x[53] & ~x[54] & ~x[56] & ~x[60];
			partial_clause[316] 	= partial_clause_prev[316] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[13] & ~x[18] & ~x[33] & ~x[36] & ~x[39] & ~x[41] & ~x[43] & ~x[46] & ~x[47] & ~x[60] & ~x[61];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[20] & ~x[26] & ~x[28] & ~x[33] & ~x[47] & ~x[63];
			partial_clause[318] 	= partial_clause_prev[318] & ~x[24] & ~x[51];
			partial_clause[319] 	= partial_clause_prev[319] & ~x[25] & ~x[37] & ~x[47] & ~x[58];
			partial_clause[320] 	= partial_clause_prev[320] & ~x[10] & ~x[14] & ~x[15] & ~x[45] & ~x[46];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[14] & ~x[21] & ~x[42] & ~x[45] & ~x[48] & ~x[49];
			partial_clause[322] 	= partial_clause_prev[322] & 1'b1;
			partial_clause[323] 	= partial_clause_prev[323] & ~x[6] & ~x[23] & ~x[27] & ~x[28];
			partial_clause[324] 	= partial_clause_prev[324] & 1'b1;
			partial_clause[325] 	= partial_clause_prev[325] & ~x[11] & ~x[13] & ~x[16] & ~x[18] & ~x[38] & ~x[41] & ~x[45] & ~x[62] & ~x[63];
			partial_clause[326] 	= partial_clause_prev[326] & ~x[1] & ~x[5] & ~x[12] & ~x[13] & ~x[14] & ~x[16] & ~x[18] & ~x[37] & ~x[38] & ~x[39] & ~x[41];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[34] & ~x[39] & ~x[43] & ~x[59];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[18] & ~x[38] & ~x[40] & ~x[45];
			partial_clause[329] 	= partial_clause_prev[329] & ~x[56];
			partial_clause[330] 	= partial_clause_prev[330] & ~x[41];
			partial_clause[331] 	= partial_clause_prev[331] & ~x[9] & ~x[15] & ~x[36] & ~x[39];
			partial_clause[332] 	= partial_clause_prev[332] & ~x[11] & ~x[63];
			partial_clause[333] 	= partial_clause_prev[333] & 1'b1;
			partial_clause[334] 	= partial_clause_prev[334] & ~x[12] & ~x[45];
			partial_clause[335] 	= partial_clause_prev[335] & ~x[5] & ~x[17] & ~x[36] & ~x[63];
			partial_clause[336] 	= partial_clause_prev[336] & 1'b1;
			partial_clause[337] 	= partial_clause_prev[337] & ~x[6] & ~x[16] & ~x[39] & ~x[40] & ~x[45];
			partial_clause[338] 	= partial_clause_prev[338] & 1'b1;
			partial_clause[339] 	= partial_clause_prev[339] & ~x[11] & ~x[12] & ~x[13] & ~x[16] & ~x[17] & ~x[18] & ~x[20] & ~x[21] & ~x[38] & ~x[40] & ~x[42] & ~x[44] & ~x[45] & ~x[48];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[0] & ~x[1] & ~x[2] & ~x[6] & ~x[13] & ~x[15] & ~x[20] & ~x[26] & ~x[27] & ~x[28] & ~x[30] & ~x[34] & ~x[39] & ~x[46] & ~x[47];
			partial_clause[341] 	= partial_clause_prev[341] & x[54];
			partial_clause[342] 	= partial_clause_prev[342] & ~x[11] & ~x[14] & ~x[17] & ~x[38] & ~x[45] & x[56];
			partial_clause[343] 	= partial_clause_prev[343] & ~x[5] & ~x[6] & ~x[35] & ~x[36] & ~x[39] & ~x[41];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[9] & ~x[23];
			partial_clause[345] 	= partial_clause_prev[345] & ~x[1] & ~x[31];
			partial_clause[346] 	= partial_clause_prev[346] & ~x[1] & ~x[32];
			partial_clause[347] 	= partial_clause_prev[347] & ~x[9] & ~x[12] & ~x[18];
			partial_clause[348] 	= partial_clause_prev[348] & ~x[7] & ~x[8] & ~x[12] & ~x[15] & ~x[40];
			partial_clause[349] 	= partial_clause_prev[349] & ~x[1] & ~x[12] & ~x[28] & ~x[32];
			partial_clause[350] 	= partial_clause_prev[350] & ~x[1] & ~x[4] & ~x[6] & ~x[7] & ~x[10] & ~x[11] & ~x[13] & ~x[16] & ~x[17] & ~x[34] & ~x[36] & ~x[37] & ~x[40] & ~x[44] & ~x[46] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[351] 	= partial_clause_prev[351] & 1'b1;
			partial_clause[352] 	= partial_clause_prev[352] & ~x[19];
			partial_clause[353] 	= partial_clause_prev[353] & ~x[19] & ~x[26];
			partial_clause[354] 	= partial_clause_prev[354] & ~x[8] & ~x[14] & ~x[17] & ~x[35] & ~x[40] & ~x[45];
			partial_clause[355] 	= partial_clause_prev[355] & ~x[2] & ~x[31] & ~x[35];
			partial_clause[356] 	= partial_clause_prev[356] & 1'b1;
			partial_clause[357] 	= partial_clause_prev[357] & 1'b1;
			partial_clause[358] 	= partial_clause_prev[358] & ~x[4] & ~x[5] & ~x[9] & ~x[10] & ~x[12] & ~x[47];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[3] & ~x[5] & ~x[8] & ~x[37] & ~x[38];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[0] & ~x[2] & ~x[13] & ~x[16] & ~x[18] & ~x[19] & ~x[21] & ~x[23] & ~x[25] & ~x[26] & ~x[32] & ~x[44] & ~x[59] & ~x[61];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[18] & ~x[44] & ~x[46];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[1] & ~x[5] & ~x[19] & ~x[42] & ~x[47];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[4] & ~x[13] & ~x[31] & ~x[32] & ~x[35] & ~x[41] & ~x[47];
			partial_clause[364] 	= partial_clause_prev[364] & ~x[23] & ~x[44];
			partial_clause[365] 	= partial_clause_prev[365] & 1'b1;
			partial_clause[366] 	= partial_clause_prev[366] & ~x[0] & ~x[3] & ~x[13] & ~x[20] & ~x[21] & ~x[29] & ~x[37] & ~x[38] & ~x[40] & ~x[42];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[10] & ~x[13] & ~x[38] & ~x[40] & ~x[44] & ~x[51];
			partial_clause[368] 	= partial_clause_prev[368] & ~x[60];
			partial_clause[369] 	= partial_clause_prev[369] & ~x[11] & ~x[12] & ~x[14] & ~x[15] & ~x[19] & ~x[22] & ~x[37];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[21] & ~x[23] & ~x[36] & ~x[39] & ~x[49] & ~x[62] & ~x[63];
			partial_clause[371] 	= partial_clause_prev[371] & ~x[42];
			partial_clause[372] 	= partial_clause_prev[372] & ~x[5] & ~x[12] & ~x[30] & ~x[34];
			partial_clause[373] 	= partial_clause_prev[373] & ~x[49] & ~x[56];
			partial_clause[374] 	= partial_clause_prev[374] & ~x[9] & ~x[40];
			partial_clause[375] 	= partial_clause_prev[375] & ~x[1];
			partial_clause[376] 	= partial_clause_prev[376] & ~x[3] & ~x[4] & ~x[8] & ~x[9] & ~x[11] & ~x[35] & ~x[63];
			partial_clause[377] 	= partial_clause_prev[377] & ~x[7] & ~x[8] & ~x[39];
			partial_clause[378] 	= partial_clause_prev[378] & ~x[13];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[42];
			partial_clause[380] 	= partial_clause_prev[380] & ~x[57];
			partial_clause[381] 	= partial_clause_prev[381] & ~x[3] & ~x[6] & ~x[8] & ~x[10] & ~x[16] & ~x[39] & ~x[40] & ~x[41] & ~x[42];
			partial_clause[382] 	= partial_clause_prev[382] & 1'b1;
			partial_clause[383] 	= partial_clause_prev[383] & 1'b1;
			partial_clause[384] 	= partial_clause_prev[384] & 1'b1;
			partial_clause[385] 	= partial_clause_prev[385] & x[25] & x[26] & x[27] & ~x[32] & ~x[33];
			partial_clause[386] 	= partial_clause_prev[386] & ~x[6];
			partial_clause[387] 	= partial_clause_prev[387] & ~x[8] & ~x[11] & ~x[14] & ~x[15] & ~x[17] & ~x[35] & ~x[42];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[13] & ~x[16] & ~x[17] & ~x[19] & ~x[20] & ~x[38] & ~x[40] & ~x[41] & ~x[43] & ~x[46];
			partial_clause[389] 	= partial_clause_prev[389] & ~x[53];
			partial_clause[390] 	= partial_clause_prev[390] & ~x[7] & ~x[15] & ~x[17] & ~x[33] & ~x[35] & ~x[36] & ~x[45] & ~x[46] & x[53];
			partial_clause[391] 	= partial_clause_prev[391] & ~x[54];
			partial_clause[392] 	= partial_clause_prev[392] & 1'b1;
			partial_clause[393] 	= partial_clause_prev[393] & 1'b1;
			partial_clause[394] 	= partial_clause_prev[394] & ~x[60];
			partial_clause[395] 	= partial_clause_prev[395] & 1'b1;
			partial_clause[396] 	= partial_clause_prev[396] & 1'b1;
			partial_clause[397] 	= partial_clause_prev[397] & ~x[23];
			partial_clause[398] 	= partial_clause_prev[398] & 1'b1;
			partial_clause[399] 	= partial_clause_prev[399] & ~x[60];
			partial_clause[400] 	= partial_clause_prev[400] & ~x[9] & ~x[18] & ~x[33] & ~x[43] & ~x[48];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[10] & ~x[14] & ~x[15] & ~x[38] & ~x[40];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[10] & ~x[11] & ~x[12] & ~x[18] & ~x[21] & ~x[37] & ~x[38];
			partial_clause[403] 	= partial_clause_prev[403] & ~x[8];
			partial_clause[404] 	= partial_clause_prev[404] & 1'b1;
			partial_clause[405] 	= partial_clause_prev[405] & ~x[24] & ~x[40] & ~x[41] & ~x[50];
			partial_clause[406] 	= partial_clause_prev[406] & ~x[9] & ~x[41] & ~x[48];
			partial_clause[407] 	= partial_clause_prev[407] & ~x[17];
			partial_clause[408] 	= partial_clause_prev[408] & 1'b1;
			partial_clause[409] 	= partial_clause_prev[409] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[18] & ~x[20] & ~x[38] & ~x[41] & ~x[46] & ~x[47] & ~x[63];
			partial_clause[410] 	= partial_clause_prev[410] & ~x[13] & ~x[16] & ~x[18];
			partial_clause[411] 	= partial_clause_prev[411] & ~x[5] & ~x[46] & ~x[63];
			partial_clause[412] 	= partial_clause_prev[412] & ~x[10] & ~x[12] & ~x[13] & ~x[14] & ~x[16] & ~x[22] & ~x[43] & ~x[46] & ~x[48] & ~x[49];
			partial_clause[413] 	= partial_clause_prev[413] & ~x[14] & ~x[43];
			partial_clause[414] 	= partial_clause_prev[414] & ~x[3] & ~x[4] & ~x[7] & ~x[10] & ~x[11] & ~x[13] & ~x[15] & ~x[16] & ~x[23] & ~x[27] & ~x[39] & ~x[42] & ~x[43] & ~x[47] & ~x[48] & ~x[50];
			partial_clause[415] 	= partial_clause_prev[415] & ~x[11] & ~x[16] & ~x[33] & ~x[45];
			partial_clause[416] 	= partial_clause_prev[416] & ~x[17] & ~x[18] & ~x[38] & ~x[41];
			partial_clause[417] 	= partial_clause_prev[417] & ~x[4] & ~x[16];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[7] & ~x[14] & ~x[19] & ~x[28] & ~x[38] & ~x[46] & ~x[62];
			partial_clause[419] 	= partial_clause_prev[419] & 1'b1;
			partial_clause[420] 	= partial_clause_prev[420] & 1'b1;
			partial_clause[421] 	= partial_clause_prev[421] & ~x[1] & ~x[5] & ~x[28] & ~x[31] & ~x[38] & ~x[39] & ~x[44];
			partial_clause[422] 	= partial_clause_prev[422] & ~x[11] & ~x[33] & ~x[34] & ~x[38];
			partial_clause[423] 	= partial_clause_prev[423] & ~x[5] & ~x[37];
			partial_clause[424] 	= partial_clause_prev[424] & ~x[25] & ~x[28] & ~x[48];
			partial_clause[425] 	= partial_clause_prev[425] & ~x[12] & ~x[36];
			partial_clause[426] 	= partial_clause_prev[426] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[12] & ~x[16] & ~x[17] & ~x[39] & ~x[42];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[7] & ~x[8] & ~x[11] & ~x[12] & ~x[20] & ~x[42];
			partial_clause[428] 	= partial_clause_prev[428] & 1'b1;
			partial_clause[429] 	= partial_clause_prev[429] & 1'b1;
			partial_clause[430] 	= partial_clause_prev[430] & ~x[4] & ~x[43] & ~x[45];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[10];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[12] & ~x[13] & ~x[15] & ~x[17] & ~x[20] & ~x[38] & ~x[44];
			partial_clause[433] 	= partial_clause_prev[433] & ~x[4];
			partial_clause[434] 	= partial_clause_prev[434] & ~x[13] & ~x[28] & ~x[33];
			partial_clause[435] 	= partial_clause_prev[435] & ~x[4] & ~x[6] & ~x[10] & ~x[12] & ~x[16] & ~x[18] & ~x[33] & ~x[37] & ~x[40] & ~x[41] & ~x[42] & ~x[45];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[6] & ~x[10] & ~x[12] & ~x[38] & ~x[63];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[16] & ~x[18] & ~x[21] & ~x[41] & ~x[43] & ~x[44] & ~x[47] & ~x[49];
			partial_clause[438] 	= partial_clause_prev[438] & ~x[16] & ~x[33];
			partial_clause[439] 	= partial_clause_prev[439] & ~x[5] & ~x[9] & ~x[15] & ~x[41];
			partial_clause[440] 	= partial_clause_prev[440] & ~x[42] & ~x[63];
			partial_clause[441] 	= partial_clause_prev[441] & ~x[18];
			partial_clause[442] 	= partial_clause_prev[442] & ~x[51];
			partial_clause[443] 	= partial_clause_prev[443] & ~x[0] & ~x[9] & ~x[15] & ~x[31] & ~x[37] & ~x[38] & ~x[41] & ~x[61];
			partial_clause[444] 	= partial_clause_prev[444] & 1'b1;
			partial_clause[445] 	= partial_clause_prev[445] & 1'b1;
			partial_clause[446] 	= partial_clause_prev[446] & ~x[11] & ~x[39] & ~x[40];
			partial_clause[447] 	= partial_clause_prev[447] & ~x[8] & ~x[11] & ~x[17] & ~x[39] & ~x[44] & ~x[47];
			partial_clause[448] 	= partial_clause_prev[448] & ~x[25] & ~x[49] & ~x[52] & ~x[55];
			partial_clause[449] 	= partial_clause_prev[449] & ~x[13] & ~x[39] & ~x[41];
			partial_clause[450] 	= partial_clause_prev[450] & ~x[9] & ~x[28] & ~x[33] & ~x[38] & ~x[39] & ~x[45];
			partial_clause[451] 	= partial_clause_prev[451] & ~x[60];
			partial_clause[452] 	= partial_clause_prev[452] & 1'b1;
			partial_clause[453] 	= partial_clause_prev[453] & ~x[0] & ~x[11] & ~x[46];
			partial_clause[454] 	= partial_clause_prev[454] & ~x[39] & ~x[53];
			partial_clause[455] 	= partial_clause_prev[455] & ~x[20] & ~x[49];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[6] & ~x[7] & ~x[39] & ~x[40] & ~x[45] & ~x[49];
			partial_clause[457] 	= partial_clause_prev[457] & 1'b1;
			partial_clause[458] 	= partial_clause_prev[458] & ~x[37] & ~x[42] & ~x[62];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[10] & ~x[19] & ~x[20] & ~x[42] & ~x[47] & ~x[50] & ~x[51];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[2] & ~x[5] & ~x[17] & ~x[18] & ~x[36] & ~x[38] & ~x[39] & ~x[41] & ~x[44] & ~x[46];
			partial_clause[461] 	= partial_clause_prev[461] & ~x[5] & ~x[39] & ~x[62];
			partial_clause[462] 	= partial_clause_prev[462] & 1'b1;
			partial_clause[463] 	= partial_clause_prev[463] & 1'b1;
			partial_clause[464] 	= partial_clause_prev[464] & ~x[7] & ~x[14];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[12] & ~x[15] & ~x[41] & ~x[42];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[5] & ~x[6] & ~x[8] & ~x[16] & ~x[19] & ~x[41] & ~x[45];
			partial_clause[467] 	= partial_clause_prev[467] & ~x[7] & ~x[9] & ~x[35];
			partial_clause[468] 	= partial_clause_prev[468] & ~x[11] & ~x[44];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[3] & ~x[8] & ~x[35] & ~x[37] & ~x[43] & ~x[45] & ~x[62];
			partial_clause[470] 	= partial_clause_prev[470] & ~x[46];
			partial_clause[471] 	= partial_clause_prev[471] & ~x[14] & ~x[16] & ~x[18] & ~x[21] & ~x[34] & ~x[38] & ~x[39] & ~x[40] & ~x[42] & ~x[49];
			partial_clause[472] 	= partial_clause_prev[472] & ~x[7] & ~x[18] & ~x[23] & ~x[24] & ~x[26] & ~x[27] & ~x[32] & ~x[62];
			partial_clause[473] 	= partial_clause_prev[473] & ~x[1] & ~x[2] & ~x[6] & ~x[10] & ~x[31] & ~x[42] & ~x[59] & ~x[60] & ~x[61] & ~x[63];
			partial_clause[474] 	= partial_clause_prev[474] & 1'b1;
			partial_clause[475] 	= partial_clause_prev[475] & ~x[28] & ~x[30] & ~x[42] & ~x[48] & ~x[62];
			partial_clause[476] 	= partial_clause_prev[476] & ~x[44] & ~x[45];
			partial_clause[477] 	= partial_clause_prev[477] & ~x[10] & ~x[13] & ~x[42];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[9] & ~x[10] & ~x[13] & ~x[15] & ~x[39];
			partial_clause[479] 	= partial_clause_prev[479] & 1'b1;
			partial_clause[480] 	= partial_clause_prev[480] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[20] & ~x[32] & ~x[33] & ~x[34] & ~x[36] & ~x[38] & ~x[39] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[45] & ~x[63];
			partial_clause[481] 	= partial_clause_prev[481] & ~x[9] & x[25];
			partial_clause[482] 	= partial_clause_prev[482] & ~x[9] & ~x[35] & ~x[36];
			partial_clause[483] 	= partial_clause_prev[483] & ~x[13];
			partial_clause[484] 	= partial_clause_prev[484] & ~x[12];
			partial_clause[485] 	= partial_clause_prev[485] & 1'b1;
			partial_clause[486] 	= partial_clause_prev[486] & ~x[10] & ~x[11] & ~x[36] & ~x[42] & ~x[43];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[9] & ~x[40] & ~x[41] & ~x[46];
			partial_clause[488] 	= partial_clause_prev[488] & ~x[53];
			partial_clause[489] 	= partial_clause_prev[489] & 1'b1;
			partial_clause[490] 	= partial_clause_prev[490] & 1'b1;
			partial_clause[491] 	= partial_clause_prev[491] & ~x[28] & ~x[42];
			partial_clause[492] 	= partial_clause_prev[492] & ~x[3] & ~x[14] & ~x[15] & ~x[16] & ~x[62];
			partial_clause[493] 	= partial_clause_prev[493] & 1'b1;
			partial_clause[494] 	= partial_clause_prev[494] & ~x[7] & ~x[35] & x[56];
			partial_clause[495] 	= partial_clause_prev[495] & ~x[3] & ~x[30] & ~x[32] & ~x[43];
			partial_clause[496] 	= partial_clause_prev[496] & ~x[25];
			partial_clause[497] 	= partial_clause_prev[497] & ~x[1];
			partial_clause[498] 	= partial_clause_prev[498] & 1'b1;
			partial_clause[499] 	= partial_clause_prev[499] & ~x[22];
		end
	end
endmodule


module HCB_3 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[2] & ~x[3] & ~x[6] & ~x[7] & ~x[32] & ~x[33] & ~x[59] & ~x[61] & ~x[63];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[0] & ~x[26] & ~x[59];
			partial_clause[2] 	= partial_clause_prev[2] & ~x[56];
			partial_clause[3] 	= partial_clause_prev[3] & ~x[11] & ~x[13] & x[18] & ~x[31];
			partial_clause[4] 	= partial_clause_prev[4] & ~x[3];
			partial_clause[5] 	= partial_clause_prev[5] & ~x[1] & ~x[6] & ~x[10] & ~x[28] & ~x[31] & ~x[33] & ~x[59];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[58] & ~x[60];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[9] & ~x[10] & ~x[28] & ~x[36] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[60];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[7] & ~x[10] & ~x[39] & x[49] & x[50] & ~x[60];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[4] & ~x[10] & ~x[32] & ~x[34] & ~x[62];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[6] & ~x[31] & ~x[36] & ~x[60];
			partial_clause[11] 	= partial_clause_prev[11] & ~x[1] & ~x[4] & ~x[10] & ~x[12] & ~x[13] & ~x[33] & ~x[35] & ~x[58];
			partial_clause[12] 	= partial_clause_prev[12] & ~x[5] & ~x[30] & ~x[36] & x[49] & ~x[56];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[0] & ~x[5] & ~x[10] & ~x[27] & ~x[35] & ~x[39];
			partial_clause[14] 	= partial_clause_prev[14] & 1'b1;
			partial_clause[15] 	= partial_clause_prev[15] & ~x[7];
			partial_clause[16] 	= partial_clause_prev[16] & ~x[27] & ~x[28] & ~x[61];
			partial_clause[17] 	= partial_clause_prev[17] & 1'b1;
			partial_clause[18] 	= partial_clause_prev[18] & ~x[3] & ~x[4] & ~x[30] & ~x[32] & ~x[38] & ~x[61];
			partial_clause[19] 	= partial_clause_prev[19] & ~x[2] & ~x[3] & ~x[4] & ~x[7] & ~x[31] & ~x[59];
			partial_clause[20] 	= partial_clause_prev[20] & ~x[33];
			partial_clause[21] 	= partial_clause_prev[21] & ~x[4] & ~x[37];
			partial_clause[22] 	= partial_clause_prev[22] & ~x[34];
			partial_clause[23] 	= partial_clause_prev[23] & ~x[2] & ~x[4] & ~x[5] & ~x[7] & ~x[26] & ~x[28] & ~x[31] & ~x[34] & ~x[55] & ~x[56] & ~x[58] & ~x[59] & ~x[63];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[3] & ~x[4] & ~x[5] & ~x[31] & ~x[32] & ~x[34] & ~x[35] & ~x[37] & ~x[59] & ~x[60] & ~x[63];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[4] & ~x[6] & ~x[7] & ~x[10] & ~x[12] & ~x[26] & ~x[27] & ~x[31] & ~x[59] & ~x[61] & ~x[62];
			partial_clause[26] 	= partial_clause_prev[26] & x[20] & x[22];
			partial_clause[27] 	= partial_clause_prev[27] & ~x[1] & ~x[8] & ~x[9] & ~x[22] & ~x[48] & ~x[59] & ~x[60];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[3] & ~x[10] & ~x[15] & ~x[35] & ~x[39] & ~x[41];
			partial_clause[29] 	= partial_clause_prev[29] & ~x[3] & x[18] & ~x[62];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[6];
			partial_clause[31] 	= partial_clause_prev[31] & ~x[34] & ~x[36];
			partial_clause[32] 	= partial_clause_prev[32] & ~x[4] & ~x[5] & ~x[34] & ~x[35];
			partial_clause[33] 	= partial_clause_prev[33] & x[46];
			partial_clause[34] 	= partial_clause_prev[34] & ~x[2] & ~x[5] & ~x[8] & x[17] & x[18] & ~x[27] & ~x[29] & ~x[33] & ~x[35] & ~x[52] & ~x[54] & ~x[55] & ~x[57] & ~x[59];
			partial_clause[35] 	= partial_clause_prev[35] & x[18] & ~x[63];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[3] & ~x[4] & ~x[60];
			partial_clause[37] 	= partial_clause_prev[37] & ~x[27];
			partial_clause[38] 	= partial_clause_prev[38] & ~x[7] & ~x[10] & ~x[33] & ~x[36] & ~x[59] & ~x[62] & ~x[63];
			partial_clause[39] 	= partial_clause_prev[39] & ~x[56] & ~x[58];
			partial_clause[40] 	= partial_clause_prev[40] & ~x[30] & ~x[34] & ~x[62];
			partial_clause[41] 	= partial_clause_prev[41] & 1'b1;
			partial_clause[42] 	= partial_clause_prev[42] & ~x[5];
			partial_clause[43] 	= partial_clause_prev[43] & 1'b1;
			partial_clause[44] 	= partial_clause_prev[44] & 1'b1;
			partial_clause[45] 	= partial_clause_prev[45] & ~x[7] & ~x[55];
			partial_clause[46] 	= partial_clause_prev[46] & ~x[0] & ~x[27] & ~x[28] & ~x[56] & ~x[59];
			partial_clause[47] 	= partial_clause_prev[47] & 1'b1;
			partial_clause[48] 	= partial_clause_prev[48] & 1'b1;
			partial_clause[49] 	= partial_clause_prev[49] & ~x[47] & x[50] & ~x[63];
			partial_clause[50] 	= partial_clause_prev[50] & ~x[61];
			partial_clause[51] 	= partial_clause_prev[51] & 1'b1;
			partial_clause[52] 	= partial_clause_prev[52] & 1'b1;
			partial_clause[53] 	= partial_clause_prev[53] & ~x[11];
			partial_clause[54] 	= partial_clause_prev[54] & ~x[58];
			partial_clause[55] 	= partial_clause_prev[55] & 1'b1;
			partial_clause[56] 	= partial_clause_prev[56] & ~x[19] & ~x[47];
			partial_clause[57] 	= partial_clause_prev[57] & ~x[29] & ~x[32] & ~x[33] & ~x[35] & ~x[52] & ~x[55] & ~x[57] & ~x[58] & ~x[61];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[10] & ~x[12];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[32] & ~x[62];
			partial_clause[60] 	= partial_clause_prev[60] & ~x[3];
			partial_clause[61] 	= partial_clause_prev[61] & ~x[11] & ~x[55] & ~x[59];
			partial_clause[62] 	= partial_clause_prev[62] & ~x[11] & ~x[29] & ~x[55] & ~x[56];
			partial_clause[63] 	= partial_clause_prev[63] & 1'b1;
			partial_clause[64] 	= partial_clause_prev[64] & x[43] & x[47];
			partial_clause[65] 	= partial_clause_prev[65] & ~x[25];
			partial_clause[66] 	= partial_clause_prev[66] & 1'b1;
			partial_clause[67] 	= partial_clause_prev[67] & 1'b1;
			partial_clause[68] 	= partial_clause_prev[68] & ~x[35];
			partial_clause[69] 	= partial_clause_prev[69] & ~x[4] & ~x[8] & ~x[26] & ~x[33] & ~x[36];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[1] & ~x[2] & ~x[7] & ~x[9] & ~x[14] & ~x[30] & ~x[40];
			partial_clause[71] 	= partial_clause_prev[71] & ~x[33];
			partial_clause[72] 	= partial_clause_prev[72] & ~x[1] & x[52] & ~x[56];
			partial_clause[73] 	= partial_clause_prev[73] & ~x[16];
			partial_clause[74] 	= partial_clause_prev[74] & ~x[3] & ~x[31] & ~x[33] & ~x[56];
			partial_clause[75] 	= partial_clause_prev[75] & ~x[4] & ~x[9] & ~x[12] & ~x[15] & ~x[39] & ~x[41];
			partial_clause[76] 	= partial_clause_prev[76] & ~x[1] & ~x[6] & ~x[30] & ~x[31] & ~x[33] & ~x[63];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[51] & ~x[53];
			partial_clause[78] 	= partial_clause_prev[78] & 1'b1;
			partial_clause[79] 	= partial_clause_prev[79] & ~x[1] & ~x[5] & ~x[26] & ~x[33];
			partial_clause[80] 	= partial_clause_prev[80] & ~x[20] & ~x[21] & ~x[48] & ~x[49];
			partial_clause[81] 	= partial_clause_prev[81] & 1'b1;
			partial_clause[82] 	= partial_clause_prev[82] & 1'b1;
			partial_clause[83] 	= partial_clause_prev[83] & 1'b1;
			partial_clause[84] 	= partial_clause_prev[84] & ~x[2] & x[44] & x[46] & ~x[62];
			partial_clause[85] 	= partial_clause_prev[85] & x[16] & ~x[31] & ~x[57] & ~x[58];
			partial_clause[86] 	= partial_clause_prev[86] & ~x[2] & ~x[5] & ~x[31] & ~x[36];
			partial_clause[87] 	= partial_clause_prev[87] & ~x[9] & ~x[31] & ~x[38] & ~x[53] & ~x[62];
			partial_clause[88] 	= partial_clause_prev[88] & ~x[4] & ~x[8] & x[22] & ~x[29] & ~x[35] & ~x[62];
			partial_clause[89] 	= partial_clause_prev[89] & ~x[63];
			partial_clause[90] 	= partial_clause_prev[90] & ~x[19];
			partial_clause[91] 	= partial_clause_prev[91] & x[22] & ~x[33] & x[51];
			partial_clause[92] 	= partial_clause_prev[92] & ~x[38] & ~x[41] & x[48] & ~x[60] & ~x[63];
			partial_clause[93] 	= partial_clause_prev[93] & ~x[0] & ~x[2] & ~x[4] & ~x[6] & ~x[10] & ~x[29] & ~x[31] & ~x[32] & ~x[35] & ~x[54] & ~x[58] & ~x[59];
			partial_clause[94] 	= partial_clause_prev[94] & 1'b1;
			partial_clause[95] 	= partial_clause_prev[95] & ~x[7] & ~x[35] & ~x[41] & ~x[56] & ~x[58];
			partial_clause[96] 	= partial_clause_prev[96] & 1'b1;
			partial_clause[97] 	= partial_clause_prev[97] & ~x[3] & ~x[6] & ~x[7] & ~x[9] & ~x[33] & ~x[36] & ~x[58];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[1] & ~x[5] & ~x[8] & ~x[31] & ~x[34] & ~x[36];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[1] & ~x[3] & ~x[4] & ~x[6] & ~x[28] & ~x[29] & ~x[31] & ~x[56] & ~x[57] & ~x[63];
			partial_clause[100] 	= partial_clause_prev[100] & ~x[39] & ~x[59];
			partial_clause[101] 	= partial_clause_prev[101] & 1'b1;
			partial_clause[102] 	= partial_clause_prev[102] & ~x[55];
			partial_clause[103] 	= partial_clause_prev[103] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[7] & ~x[8] & ~x[9] & ~x[12] & ~x[29] & ~x[31] & ~x[32] & ~x[34] & ~x[39];
			partial_clause[104] 	= partial_clause_prev[104] & ~x[7] & ~x[10] & ~x[38];
			partial_clause[105] 	= partial_clause_prev[105] & ~x[0] & ~x[1] & ~x[26] & ~x[29] & ~x[34] & ~x[37] & ~x[38] & ~x[55];
			partial_clause[106] 	= partial_clause_prev[106] & ~x[1] & ~x[48] & ~x[55];
			partial_clause[107] 	= partial_clause_prev[107] & ~x[7] & ~x[58] & ~x[61];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[3] & ~x[26] & ~x[28] & ~x[29] & ~x[33] & ~x[35] & ~x[58] & ~x[61] & ~x[63];
			partial_clause[109] 	= partial_clause_prev[109] & ~x[46];
			partial_clause[110] 	= partial_clause_prev[110] & ~x[24] & ~x[27];
			partial_clause[111] 	= partial_clause_prev[111] & 1'b1;
			partial_clause[112] 	= partial_clause_prev[112] & ~x[52] & ~x[59];
			partial_clause[113] 	= partial_clause_prev[113] & ~x[31];
			partial_clause[114] 	= partial_clause_prev[114] & 1'b1;
			partial_clause[115] 	= partial_clause_prev[115] & ~x[1] & ~x[2] & ~x[3] & ~x[33] & ~x[55] & ~x[57] & ~x[58];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[0] & ~x[1] & ~x[4] & ~x[5] & ~x[7] & x[20] & ~x[37] & ~x[40];
			partial_clause[117] 	= partial_clause_prev[117] & ~x[44];
			partial_clause[118] 	= partial_clause_prev[118] & ~x[3] & ~x[8] & ~x[59];
			partial_clause[119] 	= partial_clause_prev[119] & ~x[1] & ~x[2] & ~x[8] & ~x[11] & ~x[31] & ~x[38] & ~x[40];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[3] & ~x[4] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[30] & ~x[31] & ~x[32] & ~x[34] & ~x[36] & ~x[60] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[3] & ~x[31] & ~x[60] & ~x[63];
			partial_clause[122] 	= partial_clause_prev[122] & ~x[35] & ~x[43];
			partial_clause[123] 	= partial_clause_prev[123] & ~x[2] & ~x[29] & ~x[30] & ~x[31] & ~x[61];
			partial_clause[124] 	= partial_clause_prev[124] & 1'b1;
			partial_clause[125] 	= partial_clause_prev[125] & ~x[8] & ~x[34];
			partial_clause[126] 	= partial_clause_prev[126] & ~x[1] & ~x[51];
			partial_clause[127] 	= partial_clause_prev[127] & ~x[0] & ~x[1] & ~x[4] & ~x[8] & ~x[9] & ~x[27] & ~x[30] & ~x[31] & ~x[33] & ~x[56] & ~x[61] & ~x[62];
			partial_clause[128] 	= partial_clause_prev[128] & ~x[25] & ~x[36] & x[43] & ~x[54] & ~x[56] & ~x[58] & ~x[61];
			partial_clause[129] 	= partial_clause_prev[129] & ~x[1] & ~x[4] & ~x[6] & ~x[10] & ~x[28];
			partial_clause[130] 	= partial_clause_prev[130] & ~x[0] & ~x[26] & ~x[27] & ~x[34] & ~x[57];
			partial_clause[131] 	= partial_clause_prev[131] & 1'b1;
			partial_clause[132] 	= partial_clause_prev[132] & ~x[3] & ~x[4] & ~x[10] & ~x[22] & ~x[23] & ~x[33] & ~x[38] & ~x[51];
			partial_clause[133] 	= partial_clause_prev[133] & ~x[3] & ~x[4] & ~x[31];
			partial_clause[134] 	= partial_clause_prev[134] & ~x[1] & ~x[2] & ~x[3] & ~x[5] & ~x[6] & ~x[31] & ~x[34] & ~x[37] & ~x[59] & ~x[62];
			partial_clause[135] 	= partial_clause_prev[135] & ~x[12] & ~x[33] & ~x[34] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[136] 	= partial_clause_prev[136] & ~x[0] & ~x[1] & ~x[9] & ~x[27] & ~x[29] & ~x[30] & ~x[32] & ~x[58];
			partial_clause[137] 	= partial_clause_prev[137] & ~x[4];
			partial_clause[138] 	= partial_clause_prev[138] & ~x[33] & ~x[63];
			partial_clause[139] 	= partial_clause_prev[139] & ~x[5] & ~x[6] & ~x[23] & ~x[25] & ~x[26] & ~x[33] & ~x[53] & ~x[54] & ~x[59] & ~x[61] & ~x[62];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[4] & ~x[7] & ~x[8] & ~x[10] & ~x[11] & ~x[36] & ~x[41] & ~x[54] & ~x[55] & ~x[60];
			partial_clause[141] 	= partial_clause_prev[141] & ~x[35] & ~x[59];
			partial_clause[142] 	= partial_clause_prev[142] & ~x[4] & ~x[5] & ~x[28] & ~x[31] & ~x[34] & ~x[63];
			partial_clause[143] 	= partial_clause_prev[143] & 1'b1;
			partial_clause[144] 	= partial_clause_prev[144] & ~x[37];
			partial_clause[145] 	= partial_clause_prev[145] & 1'b1;
			partial_clause[146] 	= partial_clause_prev[146] & ~x[10] & ~x[35] & ~x[38] & ~x[60];
			partial_clause[147] 	= partial_clause_prev[147] & ~x[2] & ~x[5] & ~x[23] & ~x[29] & ~x[31] & ~x[41] & ~x[42] & ~x[52] & ~x[59];
			partial_clause[148] 	= partial_clause_prev[148] & ~x[30] & ~x[33];
			partial_clause[149] 	= partial_clause_prev[149] & ~x[59];
			partial_clause[150] 	= partial_clause_prev[150] & ~x[38] & ~x[60];
			partial_clause[151] 	= partial_clause_prev[151] & 1'b1;
			partial_clause[152] 	= partial_clause_prev[152] & 1'b1;
			partial_clause[153] 	= partial_clause_prev[153] & ~x[3] & ~x[4] & ~x[5] & ~x[26] & ~x[29] & ~x[34] & ~x[35] & ~x[57] & ~x[60];
			partial_clause[154] 	= partial_clause_prev[154] & 1'b1;
			partial_clause[155] 	= partial_clause_prev[155] & x[55];
			partial_clause[156] 	= partial_clause_prev[156] & ~x[1];
			partial_clause[157] 	= partial_clause_prev[157] & 1'b1;
			partial_clause[158] 	= partial_clause_prev[158] & ~x[3] & ~x[11] & ~x[13] & ~x[14] & ~x[33] & ~x[38] & ~x[61];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[0] & ~x[2] & ~x[3] & ~x[6] & ~x[9] & ~x[31] & ~x[35] & ~x[61] & ~x[62];
			partial_clause[160] 	= partial_clause_prev[160] & ~x[14] & ~x[33] & ~x[37] & ~x[41] & ~x[63];
			partial_clause[161] 	= partial_clause_prev[161] & ~x[1] & ~x[7] & ~x[9] & ~x[10] & ~x[28] & ~x[58];
			partial_clause[162] 	= partial_clause_prev[162] & ~x[0] & ~x[1] & ~x[8] & ~x[9] & ~x[35] & ~x[57];
			partial_clause[163] 	= partial_clause_prev[163] & 1'b1;
			partial_clause[164] 	= partial_clause_prev[164] & ~x[8] & ~x[14] & ~x[39];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[6] & ~x[7] & ~x[29];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[6] & ~x[9] & ~x[28] & ~x[32] & ~x[56] & ~x[58] & ~x[59] & ~x[63];
			partial_clause[167] 	= partial_clause_prev[167] & ~x[58];
			partial_clause[168] 	= partial_clause_prev[168] & ~x[2] & ~x[4] & ~x[33] & ~x[34];
			partial_clause[169] 	= partial_clause_prev[169] & ~x[38];
			partial_clause[170] 	= partial_clause_prev[170] & ~x[44];
			partial_clause[171] 	= partial_clause_prev[171] & ~x[7] & ~x[9] & ~x[60];
			partial_clause[172] 	= partial_clause_prev[172] & ~x[17] & ~x[44];
			partial_clause[173] 	= partial_clause_prev[173] & ~x[1] & ~x[3] & ~x[6] & ~x[31] & ~x[36] & ~x[38] & ~x[57] & ~x[62];
			partial_clause[174] 	= partial_clause_prev[174] & ~x[6];
			partial_clause[175] 	= partial_clause_prev[175] & ~x[47];
			partial_clause[176] 	= partial_clause_prev[176] & ~x[27];
			partial_clause[177] 	= partial_clause_prev[177] & ~x[0] & x[18] & x[19] & ~x[55] & ~x[62];
			partial_clause[178] 	= partial_clause_prev[178] & ~x[5] & x[20];
			partial_clause[179] 	= partial_clause_prev[179] & 1'b1;
			partial_clause[180] 	= partial_clause_prev[180] & ~x[29] & ~x[35];
			partial_clause[181] 	= partial_clause_prev[181] & 1'b1;
			partial_clause[182] 	= partial_clause_prev[182] & ~x[56];
			partial_clause[183] 	= partial_clause_prev[183] & ~x[4] & ~x[8] & ~x[9] & ~x[12] & ~x[14] & ~x[32] & ~x[35] & ~x[41] & ~x[60];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[3] & ~x[33] & ~x[36] & ~x[39] & ~x[42] & ~x[61];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[1] & ~x[3] & ~x[7] & ~x[30] & ~x[62] & ~x[63];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[1] & ~x[6] & ~x[7] & ~x[8] & ~x[10] & ~x[25] & ~x[26] & ~x[30] & ~x[52] & ~x[55] & ~x[57] & ~x[58] & ~x[63];
			partial_clause[187] 	= partial_clause_prev[187] & ~x[3] & ~x[9] & ~x[24] & ~x[26] & ~x[31] & ~x[34] & ~x[54] & ~x[58] & ~x[61];
			partial_clause[188] 	= partial_clause_prev[188] & ~x[60];
			partial_clause[189] 	= partial_clause_prev[189] & 1'b1;
			partial_clause[190] 	= partial_clause_prev[190] & ~x[1] & ~x[4] & ~x[13];
			partial_clause[191] 	= partial_clause_prev[191] & ~x[8] & ~x[32] & ~x[44] & ~x[55] & ~x[58] & ~x[61];
			partial_clause[192] 	= partial_clause_prev[192] & 1'b1;
			partial_clause[193] 	= partial_clause_prev[193] & ~x[22] & ~x[34] & ~x[51] & ~x[52] & ~x[60] & ~x[62];
			partial_clause[194] 	= partial_clause_prev[194] & 1'b1;
			partial_clause[195] 	= partial_clause_prev[195] & ~x[0] & ~x[1] & ~x[2] & ~x[6] & ~x[8] & ~x[9] & ~x[10] & ~x[30] & ~x[31] & ~x[33] & ~x[38] & ~x[57] & ~x[62];
			partial_clause[196] 	= partial_clause_prev[196] & ~x[10] & ~x[50];
			partial_clause[197] 	= partial_clause_prev[197] & ~x[0] & ~x[2] & ~x[4] & ~x[6] & ~x[9] & ~x[27] & ~x[32] & ~x[36] & ~x[39] & ~x[40];
			partial_clause[198] 	= partial_clause_prev[198] & ~x[62];
			partial_clause[199] 	= partial_clause_prev[199] & 1'b1;
			partial_clause[200] 	= partial_clause_prev[200] & ~x[31] & ~x[56];
			partial_clause[201] 	= partial_clause_prev[201] & ~x[8] & ~x[11] & ~x[33];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[3] & ~x[7] & ~x[10] & ~x[13] & ~x[38] & ~x[39] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[59] & ~x[61] & ~x[62];
			partial_clause[203] 	= partial_clause_prev[203] & ~x[1] & ~x[29] & ~x[33] & ~x[59];
			partial_clause[204] 	= partial_clause_prev[204] & ~x[3] & ~x[7] & ~x[11] & ~x[31] & ~x[33] & ~x[34] & ~x[41] & ~x[58] & ~x[61] & ~x[62];
			partial_clause[205] 	= partial_clause_prev[205] & x[22] & x[23];
			partial_clause[206] 	= partial_clause_prev[206] & ~x[7] & ~x[32] & ~x[35] & ~x[60];
			partial_clause[207] 	= partial_clause_prev[207] & ~x[1] & ~x[6] & ~x[37] & ~x[51];
			partial_clause[208] 	= partial_clause_prev[208] & ~x[0] & ~x[4] & ~x[8] & ~x[37];
			partial_clause[209] 	= partial_clause_prev[209] & ~x[13] & ~x[43];
			partial_clause[210] 	= partial_clause_prev[210] & ~x[0] & ~x[1] & ~x[31] & ~x[37] & ~x[39] & ~x[41];
			partial_clause[211] 	= partial_clause_prev[211] & 1'b1;
			partial_clause[212] 	= partial_clause_prev[212] & ~x[25] & ~x[38];
			partial_clause[213] 	= partial_clause_prev[213] & 1'b1;
			partial_clause[214] 	= partial_clause_prev[214] & ~x[11] & ~x[56];
			partial_clause[215] 	= partial_clause_prev[215] & 1'b1;
			partial_clause[216] 	= partial_clause_prev[216] & x[19];
			partial_clause[217] 	= partial_clause_prev[217] & ~x[1] & ~x[8] & ~x[26];
			partial_clause[218] 	= partial_clause_prev[218] & 1'b1;
			partial_clause[219] 	= partial_clause_prev[219] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[54];
			partial_clause[220] 	= partial_clause_prev[220] & ~x[3] & ~x[5] & ~x[9] & ~x[12] & ~x[33] & ~x[35] & ~x[60];
			partial_clause[221] 	= partial_clause_prev[221] & 1'b1;
			partial_clause[222] 	= partial_clause_prev[222] & ~x[10] & ~x[13] & ~x[56];
			partial_clause[223] 	= partial_clause_prev[223] & ~x[62] & ~x[63];
			partial_clause[224] 	= partial_clause_prev[224] & ~x[11] & ~x[28] & ~x[30] & ~x[36] & ~x[39] & ~x[62];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[0] & ~x[10] & ~x[60];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[5] & ~x[7] & ~x[8] & ~x[10] & ~x[11] & ~x[29] & ~x[30] & ~x[34] & ~x[35] & ~x[57] & ~x[58] & ~x[62] & ~x[63];
			partial_clause[227] 	= partial_clause_prev[227] & ~x[9];
			partial_clause[228] 	= partial_clause_prev[228] & ~x[6] & ~x[9] & ~x[14] & ~x[31] & ~x[36] & ~x[40] & ~x[61];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[11] & ~x[34] & ~x[37] & ~x[56];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[2] & ~x[3] & ~x[5] & ~x[8] & ~x[30] & ~x[31] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[60] & ~x[62];
			partial_clause[231] 	= partial_clause_prev[231] & ~x[0] & ~x[2] & ~x[4] & ~x[31] & ~x[35] & ~x[63];
			partial_clause[232] 	= partial_clause_prev[232] & 1'b1;
			partial_clause[233] 	= partial_clause_prev[233] & 1'b1;
			partial_clause[234] 	= partial_clause_prev[234] & ~x[25] & ~x[35] & ~x[60];
			partial_clause[235] 	= partial_clause_prev[235] & 1'b1;
			partial_clause[236] 	= partial_clause_prev[236] & 1'b1;
			partial_clause[237] 	= partial_clause_prev[237] & x[13] & x[14];
			partial_clause[238] 	= partial_clause_prev[238] & 1'b1;
			partial_clause[239] 	= partial_clause_prev[239] & 1'b1;
			partial_clause[240] 	= partial_clause_prev[240] & ~x[1] & ~x[2] & ~x[6] & ~x[11] & ~x[13] & ~x[27] & ~x[32] & ~x[39];
			partial_clause[241] 	= partial_clause_prev[241] & 1'b1;
			partial_clause[242] 	= partial_clause_prev[242] & ~x[6] & ~x[9] & ~x[10] & ~x[11] & ~x[30] & ~x[39] & ~x[59] & ~x[60];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[1] & ~x[2] & ~x[5] & ~x[7] & ~x[55] & ~x[56];
			partial_clause[244] 	= partial_clause_prev[244] & 1'b1;
			partial_clause[245] 	= partial_clause_prev[245] & 1'b1;
			partial_clause[246] 	= partial_clause_prev[246] & ~x[6] & ~x[34] & ~x[60];
			partial_clause[247] 	= partial_clause_prev[247] & ~x[9] & ~x[12] & ~x[30] & ~x[36] & ~x[60];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[0] & ~x[1] & ~x[2] & ~x[4] & ~x[7] & ~x[28] & ~x[35] & ~x[36] & ~x[55] & ~x[56] & ~x[59] & ~x[60];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[26];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[1] & ~x[2] & ~x[4] & ~x[27] & ~x[28] & ~x[31] & ~x[57] & ~x[59] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[251] 	= partial_clause_prev[251] & ~x[1];
			partial_clause[252] 	= partial_clause_prev[252] & ~x[0] & ~x[8] & ~x[9] & ~x[23] & ~x[27] & ~x[28] & ~x[29] & ~x[33] & ~x[57] & ~x[58] & ~x[61];
			partial_clause[253] 	= partial_clause_prev[253] & ~x[24] & ~x[33] & ~x[43] & x[47] & ~x[56];
			partial_clause[254] 	= partial_clause_prev[254] & ~x[4] & ~x[8] & ~x[32] & ~x[56];
			partial_clause[255] 	= partial_clause_prev[255] & ~x[0] & ~x[4] & ~x[25] & ~x[34] & ~x[55] & ~x[56] & ~x[62];
			partial_clause[256] 	= partial_clause_prev[256] & ~x[13];
			partial_clause[257] 	= partial_clause_prev[257] & ~x[7] & ~x[10] & ~x[62] & ~x[63];
			partial_clause[258] 	= partial_clause_prev[258] & 1'b1;
			partial_clause[259] 	= partial_clause_prev[259] & 1'b1;
			partial_clause[260] 	= partial_clause_prev[260] & ~x[63];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[8] & ~x[57];
			partial_clause[262] 	= partial_clause_prev[262] & x[13] & ~x[34] & ~x[36] & ~x[59];
			partial_clause[263] 	= partial_clause_prev[263] & x[44];
			partial_clause[264] 	= partial_clause_prev[264] & ~x[10] & x[20] & ~x[27];
			partial_clause[265] 	= partial_clause_prev[265] & 1'b1;
			partial_clause[266] 	= partial_clause_prev[266] & ~x[1] & ~x[2] & ~x[7] & ~x[8] & ~x[28] & ~x[33] & ~x[55] & ~x[56];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[4] & ~x[7] & ~x[8] & ~x[9] & ~x[30] & ~x[32] & ~x[34] & ~x[58] & ~x[59] & ~x[60];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[1] & ~x[2] & ~x[8] & ~x[28] & ~x[30] & ~x[34] & ~x[35] & ~x[59] & ~x[60];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[2] & ~x[4] & ~x[8] & ~x[9] & ~x[12] & ~x[30] & ~x[31] & ~x[33] & ~x[34] & ~x[35] & ~x[37] & ~x[38] & ~x[39] & ~x[58] & ~x[60] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[270] 	= partial_clause_prev[270] & ~x[22] & ~x[24];
			partial_clause[271] 	= partial_clause_prev[271] & ~x[29];
			partial_clause[272] 	= partial_clause_prev[272] & ~x[4] & ~x[32] & ~x[60] & ~x[61];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[1] & ~x[6] & ~x[7] & ~x[9] & ~x[28] & ~x[31] & ~x[35] & ~x[57] & ~x[58] & ~x[63];
			partial_clause[274] 	= partial_clause_prev[274] & ~x[0] & ~x[3];
			partial_clause[275] 	= partial_clause_prev[275] & ~x[17] & ~x[27] & ~x[45] & ~x[54];
			partial_clause[276] 	= partial_clause_prev[276] & 1'b1;
			partial_clause[277] 	= partial_clause_prev[277] & ~x[11] & ~x[12] & ~x[37];
			partial_clause[278] 	= partial_clause_prev[278] & x[17];
			partial_clause[279] 	= partial_clause_prev[279] & ~x[3] & ~x[4] & ~x[6] & ~x[11] & ~x[12] & ~x[26] & ~x[29] & ~x[39] & ~x[53] & ~x[55] & ~x[61] & ~x[62];
			partial_clause[280] 	= partial_clause_prev[280] & 1'b1;
			partial_clause[281] 	= partial_clause_prev[281] & ~x[23] & ~x[25] & ~x[31] & ~x[50] & ~x[57];
			partial_clause[282] 	= partial_clause_prev[282] & ~x[4] & ~x[27] & ~x[28] & ~x[34] & ~x[63];
			partial_clause[283] 	= partial_clause_prev[283] & ~x[58];
			partial_clause[284] 	= partial_clause_prev[284] & ~x[34] & ~x[54];
			partial_clause[285] 	= partial_clause_prev[285] & x[39] & x[40];
			partial_clause[286] 	= partial_clause_prev[286] & 1'b1;
			partial_clause[287] 	= partial_clause_prev[287] & ~x[5] & ~x[7] & ~x[8] & ~x[31] & ~x[37] & ~x[59] & ~x[60] & ~x[61];
			partial_clause[288] 	= partial_clause_prev[288] & 1'b1;
			partial_clause[289] 	= partial_clause_prev[289] & 1'b1;
			partial_clause[290] 	= partial_clause_prev[290] & ~x[23] & ~x[32];
			partial_clause[291] 	= partial_clause_prev[291] & ~x[44] & ~x[59];
			partial_clause[292] 	= partial_clause_prev[292] & ~x[34];
			partial_clause[293] 	= partial_clause_prev[293] & ~x[58] & ~x[61];
			partial_clause[294] 	= partial_clause_prev[294] & ~x[2] & ~x[39] & ~x[58] & ~x[61];
			partial_clause[295] 	= partial_clause_prev[295] & ~x[59];
			partial_clause[296] 	= partial_clause_prev[296] & 1'b1;
			partial_clause[297] 	= partial_clause_prev[297] & ~x[11];
			partial_clause[298] 	= partial_clause_prev[298] & 1'b1;
			partial_clause[299] 	= partial_clause_prev[299] & ~x[0] & ~x[1] & x[19] & ~x[32] & ~x[34] & x[46] & ~x[55];
			partial_clause[300] 	= partial_clause_prev[300] & ~x[31] & ~x[32] & ~x[47] & ~x[59] & ~x[63];
			partial_clause[301] 	= partial_clause_prev[301] & ~x[2] & ~x[6] & ~x[10] & ~x[14] & ~x[57];
			partial_clause[302] 	= partial_clause_prev[302] & ~x[7] & ~x[46];
			partial_clause[303] 	= partial_clause_prev[303] & x[46];
			partial_clause[304] 	= partial_clause_prev[304] & ~x[6];
			partial_clause[305] 	= partial_clause_prev[305] & ~x[32];
			partial_clause[306] 	= partial_clause_prev[306] & ~x[3] & ~x[5] & ~x[29] & ~x[59] & ~x[60];
			partial_clause[307] 	= partial_clause_prev[307] & ~x[1] & ~x[6] & ~x[9] & ~x[28] & ~x[33];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[0] & ~x[4] & ~x[31] & ~x[55] & ~x[57] & ~x[60];
			partial_clause[309] 	= partial_clause_prev[309] & ~x[3] & ~x[6] & ~x[57] & ~x[60];
			partial_clause[310] 	= partial_clause_prev[310] & 1'b1;
			partial_clause[311] 	= partial_clause_prev[311] & ~x[36];
			partial_clause[312] 	= partial_clause_prev[312] & ~x[61];
			partial_clause[313] 	= partial_clause_prev[313] & ~x[1] & ~x[12] & ~x[62];
			partial_clause[314] 	= partial_clause_prev[314] & ~x[6];
			partial_clause[315] 	= partial_clause_prev[315] & ~x[57];
			partial_clause[316] 	= partial_clause_prev[316] & ~x[9] & ~x[26] & ~x[30] & ~x[31] & ~x[36] & ~x[38] & ~x[52] & ~x[58] & ~x[61];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[2];
			partial_clause[318] 	= partial_clause_prev[318] & ~x[14] & ~x[42] & ~x[59];
			partial_clause[319] 	= partial_clause_prev[319] & ~x[35];
			partial_clause[320] 	= partial_clause_prev[320] & ~x[3] & ~x[28] & ~x[37] & ~x[58];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[5] & ~x[7] & ~x[30] & ~x[33] & ~x[34] & ~x[35] & ~x[58];
			partial_clause[322] 	= partial_clause_prev[322] & ~x[4] & ~x[12];
			partial_clause[323] 	= partial_clause_prev[323] & ~x[7] & ~x[60];
			partial_clause[324] 	= partial_clause_prev[324] & 1'b1;
			partial_clause[325] 	= partial_clause_prev[325] & ~x[2] & ~x[6] & ~x[7] & ~x[11] & ~x[29] & ~x[33] & ~x[34] & ~x[37] & ~x[38] & ~x[57] & ~x[58] & ~x[59] & ~x[61];
			partial_clause[326] 	= partial_clause_prev[326] & ~x[1] & ~x[8] & ~x[29] & ~x[32] & ~x[33] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[4] & ~x[8] & ~x[27] & ~x[52] & ~x[60] & ~x[61];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[3] & ~x[56] & ~x[63];
			partial_clause[329] 	= partial_clause_prev[329] & 1'b1;
			partial_clause[330] 	= partial_clause_prev[330] & ~x[4] & ~x[30] & ~x[33];
			partial_clause[331] 	= partial_clause_prev[331] & ~x[7] & ~x[33];
			partial_clause[332] 	= partial_clause_prev[332] & ~x[9] & ~x[10] & ~x[25] & ~x[26] & ~x[30] & ~x[34] & ~x[52] & ~x[57] & ~x[59] & ~x[60];
			partial_clause[333] 	= partial_clause_prev[333] & ~x[37];
			partial_clause[334] 	= partial_clause_prev[334] & ~x[60];
			partial_clause[335] 	= partial_clause_prev[335] & x[18] & ~x[26] & ~x[32];
			partial_clause[336] 	= partial_clause_prev[336] & 1'b1;
			partial_clause[337] 	= partial_clause_prev[337] & ~x[29] & ~x[30];
			partial_clause[338] 	= partial_clause_prev[338] & ~x[9];
			partial_clause[339] 	= partial_clause_prev[339] & ~x[9] & ~x[31] & ~x[38] & ~x[58] & ~x[59];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[2] & ~x[5] & ~x[7] & ~x[28] & x[46] & x[47] & ~x[57];
			partial_clause[341] 	= partial_clause_prev[341] & 1'b1;
			partial_clause[342] 	= partial_clause_prev[342] & ~x[6] & x[19] & x[20] & ~x[29] & ~x[33] & ~x[34] & ~x[38];
			partial_clause[343] 	= partial_clause_prev[343] & ~x[6] & x[20] & ~x[31] & ~x[62];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[3] & ~x[12] & ~x[13] & ~x[14] & ~x[27] & ~x[42] & ~x[55];
			partial_clause[345] 	= partial_clause_prev[345] & ~x[1] & ~x[57];
			partial_clause[346] 	= partial_clause_prev[346] & ~x[1];
			partial_clause[347] 	= partial_clause_prev[347] & ~x[1] & ~x[4] & ~x[27] & ~x[56];
			partial_clause[348] 	= partial_clause_prev[348] & ~x[5];
			partial_clause[349] 	= partial_clause_prev[349] & ~x[4] & x[51];
			partial_clause[350] 	= partial_clause_prev[350] & ~x[2] & ~x[3] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[25] & ~x[27] & ~x[28] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[35] & ~x[54] & ~x[55] & ~x[57] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[351] 	= partial_clause_prev[351] & ~x[4];
			partial_clause[352] 	= partial_clause_prev[352] & x[22];
			partial_clause[353] 	= partial_clause_prev[353] & ~x[3];
			partial_clause[354] 	= partial_clause_prev[354] & ~x[3] & ~x[6] & ~x[7] & ~x[8] & ~x[30] & ~x[34] & ~x[37];
			partial_clause[355] 	= partial_clause_prev[355] & ~x[0] & ~x[27] & ~x[31] & ~x[35] & ~x[63];
			partial_clause[356] 	= partial_clause_prev[356] & ~x[3] & ~x[5] & ~x[10] & ~x[30] & ~x[52];
			partial_clause[357] 	= partial_clause_prev[357] & 1'b1;
			partial_clause[358] 	= partial_clause_prev[358] & ~x[0] & ~x[7] & ~x[26] & ~x[27];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[3] & ~x[4] & ~x[32];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[1] & ~x[3] & ~x[5] & ~x[6] & ~x[8] & ~x[9] & ~x[27] & ~x[28] & ~x[32] & ~x[34] & ~x[36] & ~x[55] & ~x[56] & ~x[57] & ~x[58];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[6] & ~x[36] & ~x[62];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[27] & ~x[32];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[1] & ~x[7] & ~x[9] & ~x[27] & ~x[28] & ~x[35] & ~x[57];
			partial_clause[364] 	= partial_clause_prev[364] & ~x[1] & ~x[3] & ~x[14] & ~x[41];
			partial_clause[365] 	= partial_clause_prev[365] & ~x[8] & x[16];
			partial_clause[366] 	= partial_clause_prev[366] & ~x[1] & ~x[5] & ~x[31];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[10] & ~x[24] & ~x[38] & ~x[51] & ~x[63];
			partial_clause[368] 	= partial_clause_prev[368] & ~x[21] & ~x[26] & ~x[46];
			partial_clause[369] 	= partial_clause_prev[369] & ~x[0] & ~x[29] & ~x[32] & ~x[59];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[0] & ~x[6] & ~x[7] & ~x[27] & ~x[32] & ~x[34] & ~x[58] & ~x[60];
			partial_clause[371] 	= partial_clause_prev[371] & ~x[16] & ~x[24] & ~x[25] & ~x[36] & ~x[43];
			partial_clause[372] 	= partial_clause_prev[372] & ~x[63];
			partial_clause[373] 	= partial_clause_prev[373] & ~x[48];
			partial_clause[374] 	= partial_clause_prev[374] & ~x[5] & ~x[33] & ~x[59];
			partial_clause[375] 	= partial_clause_prev[375] & 1'b1;
			partial_clause[376] 	= partial_clause_prev[376] & ~x[4] & ~x[6] & ~x[29] & ~x[57];
			partial_clause[377] 	= partial_clause_prev[377] & x[21];
			partial_clause[378] 	= partial_clause_prev[378] & ~x[9] & ~x[33];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[0] & ~x[36] & ~x[56] & ~x[61] & ~x[62];
			partial_clause[380] 	= partial_clause_prev[380] & ~x[20] & ~x[48];
			partial_clause[381] 	= partial_clause_prev[381] & ~x[0] & ~x[3] & ~x[33] & ~x[34] & ~x[35] & ~x[38] & ~x[56];
			partial_clause[382] 	= partial_clause_prev[382] & 1'b1;
			partial_clause[383] 	= partial_clause_prev[383] & 1'b1;
			partial_clause[384] 	= partial_clause_prev[384] & x[43];
			partial_clause[385] 	= partial_clause_prev[385] & ~x[46];
			partial_clause[386] 	= partial_clause_prev[386] & ~x[2];
			partial_clause[387] 	= partial_clause_prev[387] & ~x[7] & ~x[36] & ~x[58];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[34] & ~x[35] & ~x[57] & ~x[59] & ~x[60];
			partial_clause[389] 	= partial_clause_prev[389] & ~x[11] & ~x[13] & ~x[15] & x[21] & ~x[41];
			partial_clause[390] 	= partial_clause_prev[390] & ~x[1] & ~x[3] & ~x[4] & ~x[10] & ~x[36] & ~x[55] & ~x[56] & ~x[58] & ~x[59];
			partial_clause[391] 	= partial_clause_prev[391] & ~x[18] & ~x[46] & x[49];
			partial_clause[392] 	= partial_clause_prev[392] & ~x[41];
			partial_clause[393] 	= partial_clause_prev[393] & 1'b1;
			partial_clause[394] 	= partial_clause_prev[394] & ~x[1] & ~x[28] & ~x[53];
			partial_clause[395] 	= partial_clause_prev[395] & ~x[9] & ~x[37];
			partial_clause[396] 	= partial_clause_prev[396] & 1'b1;
			partial_clause[397] 	= partial_clause_prev[397] & x[42] & x[45];
			partial_clause[398] 	= partial_clause_prev[398] & 1'b1;
			partial_clause[399] 	= partial_clause_prev[399] & ~x[18] & ~x[20] & ~x[22] & ~x[24] & ~x[26] & ~x[45];
			partial_clause[400] 	= partial_clause_prev[400] & ~x[29] & ~x[31] & ~x[33] & ~x[35] & ~x[62];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[7] & ~x[11] & ~x[21] & ~x[30] & ~x[33] & ~x[38];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[3] & ~x[10] & ~x[29] & ~x[32] & ~x[34];
			partial_clause[403] 	= partial_clause_prev[403] & ~x[2] & ~x[30];
			partial_clause[404] 	= partial_clause_prev[404] & ~x[23] & ~x[27] & ~x[49] & ~x[51];
			partial_clause[405] 	= partial_clause_prev[405] & ~x[8] & ~x[11] & ~x[29] & ~x[58] & ~x[60];
			partial_clause[406] 	= partial_clause_prev[406] & ~x[7] & ~x[27] & ~x[33] & ~x[60];
			partial_clause[407] 	= partial_clause_prev[407] & ~x[31] & ~x[38] & ~x[40];
			partial_clause[408] 	= partial_clause_prev[408] & ~x[1] & x[17] & ~x[63];
			partial_clause[409] 	= partial_clause_prev[409] & ~x[0] & ~x[3] & ~x[5] & ~x[8] & ~x[10] & ~x[11] & ~x[27] & ~x[29] & ~x[31] & ~x[35] & ~x[37] & ~x[38] & ~x[39] & ~x[52] & ~x[55] & ~x[56] & ~x[57] & ~x[59];
			partial_clause[410] 	= partial_clause_prev[410] & x[48] & ~x[63];
			partial_clause[411] 	= partial_clause_prev[411] & ~x[1] & ~x[26] & ~x[34] & ~x[37] & ~x[39] & ~x[54] & ~x[55] & ~x[59] & ~x[60];
			partial_clause[412] 	= partial_clause_prev[412] & ~x[1] & ~x[7] & ~x[9] & ~x[12] & ~x[31] & ~x[32] & ~x[35] & ~x[41] & ~x[56];
			partial_clause[413] 	= partial_clause_prev[413] & ~x[8] & ~x[30] & ~x[57] & ~x[59];
			partial_clause[414] 	= partial_clause_prev[414] & ~x[3] & ~x[6] & ~x[9] & ~x[13] & ~x[31] & ~x[37] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[415] 	= partial_clause_prev[415] & ~x[6] & ~x[27] & ~x[52];
			partial_clause[416] 	= partial_clause_prev[416] & ~x[5] & ~x[8] & ~x[32] & ~x[61];
			partial_clause[417] 	= partial_clause_prev[417] & ~x[36] & ~x[56];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[0] & ~x[3] & ~x[5] & ~x[6] & ~x[7] & ~x[28] & ~x[54] & ~x[56] & ~x[59];
			partial_clause[419] 	= partial_clause_prev[419] & 1'b1;
			partial_clause[420] 	= partial_clause_prev[420] & ~x[4] & ~x[63];
			partial_clause[421] 	= partial_clause_prev[421] & x[49] & ~x[61];
			partial_clause[422] 	= partial_clause_prev[422] & ~x[27] & ~x[28] & ~x[59] & ~x[60];
			partial_clause[423] 	= partial_clause_prev[423] & ~x[59];
			partial_clause[424] 	= partial_clause_prev[424] & ~x[13] & ~x[14] & ~x[58];
			partial_clause[425] 	= partial_clause_prev[425] & ~x[9] & ~x[33] & ~x[35];
			partial_clause[426] 	= partial_clause_prev[426] & ~x[4] & ~x[5] & ~x[6] & ~x[8] & ~x[35] & ~x[62] & ~x[63];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[4] & ~x[8] & ~x[32] & ~x[36] & ~x[60] & ~x[61];
			partial_clause[428] 	= partial_clause_prev[428] & ~x[30];
			partial_clause[429] 	= partial_clause_prev[429] & 1'b1;
			partial_clause[430] 	= partial_clause_prev[430] & ~x[0] & ~x[2] & ~x[9] & ~x[12] & ~x[31] & ~x[33] & ~x[39] & ~x[53] & ~x[56] & ~x[61];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[27] & ~x[60];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[0] & ~x[3] & ~x[7] & x[22] & x[23] & ~x[61] & ~x[62];
			partial_clause[433] 	= partial_clause_prev[433] & 1'b1;
			partial_clause[434] 	= partial_clause_prev[434] & ~x[32];
			partial_clause[435] 	= partial_clause_prev[435] & ~x[10] & ~x[30] & ~x[31] & ~x[32] & ~x[39] & ~x[56] & ~x[58] & ~x[59] & ~x[61] & ~x[63];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[4] & ~x[28] & ~x[56];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[5] & ~x[7] & ~x[8] & ~x[10] & ~x[12] & ~x[35] & ~x[39] & ~x[59] & ~x[60] & ~x[62];
			partial_clause[438] 	= partial_clause_prev[438] & x[20];
			partial_clause[439] 	= partial_clause_prev[439] & ~x[5] & ~x[61] & ~x[63];
			partial_clause[440] 	= partial_clause_prev[440] & ~x[59];
			partial_clause[441] 	= partial_clause_prev[441] & ~x[58] & ~x[60];
			partial_clause[442] 	= partial_clause_prev[442] & 1'b1;
			partial_clause[443] 	= partial_clause_prev[443] & ~x[1] & ~x[2] & ~x[4] & ~x[5] & ~x[7] & ~x[28] & ~x[29] & ~x[32] & ~x[57] & ~x[59];
			partial_clause[444] 	= partial_clause_prev[444] & 1'b1;
			partial_clause[445] 	= partial_clause_prev[445] & 1'b1;
			partial_clause[446] 	= partial_clause_prev[446] & ~x[34] & ~x[35] & ~x[60];
			partial_clause[447] 	= partial_clause_prev[447] & ~x[36] & ~x[63];
			partial_clause[448] 	= partial_clause_prev[448] & 1'b1;
			partial_clause[449] 	= partial_clause_prev[449] & ~x[5] & ~x[33];
			partial_clause[450] 	= partial_clause_prev[450] & ~x[10] & ~x[60] & ~x[63];
			partial_clause[451] 	= partial_clause_prev[451] & ~x[52];
			partial_clause[452] 	= partial_clause_prev[452] & 1'b1;
			partial_clause[453] 	= partial_clause_prev[453] & ~x[23] & ~x[24] & ~x[29] & ~x[31];
			partial_clause[454] 	= partial_clause_prev[454] & x[22] & ~x[63];
			partial_clause[455] 	= partial_clause_prev[455] & ~x[2] & ~x[12] & ~x[34] & ~x[36] & ~x[40] & ~x[58];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[6] & ~x[9] & ~x[10] & ~x[38] & ~x[39] & ~x[40] & ~x[57] & ~x[58] & ~x[60];
			partial_clause[457] 	= partial_clause_prev[457] & ~x[3] & ~x[33];
			partial_clause[458] 	= partial_clause_prev[458] & ~x[27] & ~x[30] & ~x[31] & ~x[37] & ~x[56] & ~x[59] & ~x[63];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[6] & ~x[14] & ~x[25] & ~x[39] & ~x[41] & ~x[42] & ~x[43] & ~x[58] & ~x[59] & ~x[60] & ~x[61];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[3] & ~x[8] & ~x[61];
			partial_clause[461] 	= partial_clause_prev[461] & x[18] & ~x[29];
			partial_clause[462] 	= partial_clause_prev[462] & ~x[32] & ~x[33];
			partial_clause[463] 	= partial_clause_prev[463] & 1'b1;
			partial_clause[464] 	= partial_clause_prev[464] & ~x[12] & ~x[30] & ~x[31] & ~x[34];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[1] & ~x[7] & ~x[32];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[0] & ~x[7] & ~x[29] & ~x[31] & ~x[33] & ~x[60] & ~x[63];
			partial_clause[467] 	= partial_clause_prev[467] & 1'b1;
			partial_clause[468] 	= partial_clause_prev[468] & ~x[8] & ~x[9] & x[20] & ~x[62];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[2] & ~x[33];
			partial_clause[470] 	= partial_clause_prev[470] & 1'b1;
			partial_clause[471] 	= partial_clause_prev[471] & ~x[8] & ~x[10] & ~x[55] & ~x[63];
			partial_clause[472] 	= partial_clause_prev[472] & ~x[34];
			partial_clause[473] 	= partial_clause_prev[473] & ~x[4] & ~x[7] & x[19] & ~x[24] & ~x[25] & ~x[26] & ~x[31] & ~x[33] & ~x[60];
			partial_clause[474] 	= partial_clause_prev[474] & ~x[63];
			partial_clause[475] 	= partial_clause_prev[475] & ~x[2] & ~x[35] & x[48] & ~x[61];
			partial_clause[476] 	= partial_clause_prev[476] & ~x[36] & ~x[59];
			partial_clause[477] 	= partial_clause_prev[477] & ~x[4] & ~x[6] & ~x[7] & ~x[28] & ~x[63];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[4] & ~x[7] & ~x[8] & ~x[17] & ~x[30] & ~x[32] & ~x[34] & ~x[36] & ~x[59];
			partial_clause[479] 	= partial_clause_prev[479] & ~x[54];
			partial_clause[480] 	= partial_clause_prev[480] & ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[7] & ~x[8] & ~x[26] & ~x[28] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[35] & ~x[54] & ~x[56] & ~x[57] & ~x[58] & ~x[59] & ~x[60] & ~x[61];
			partial_clause[481] 	= partial_clause_prev[481] & ~x[33] & ~x[34] & ~x[63];
			partial_clause[482] 	= partial_clause_prev[482] & ~x[6] & ~x[7] & ~x[32] & ~x[35];
			partial_clause[483] 	= partial_clause_prev[483] & ~x[38];
			partial_clause[484] 	= partial_clause_prev[484] & ~x[15] & ~x[52] & ~x[61] & ~x[63];
			partial_clause[485] 	= partial_clause_prev[485] & 1'b1;
			partial_clause[486] 	= partial_clause_prev[486] & ~x[5] & ~x[8] & ~x[31] & ~x[36] & ~x[60];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[8] & ~x[9] & ~x[47];
			partial_clause[488] 	= partial_clause_prev[488] & ~x[17];
			partial_clause[489] 	= partial_clause_prev[489] & ~x[29];
			partial_clause[490] 	= partial_clause_prev[490] & ~x[43];
			partial_clause[491] 	= partial_clause_prev[491] & ~x[0] & ~x[61];
			partial_clause[492] 	= partial_clause_prev[492] & ~x[26] & ~x[55];
			partial_clause[493] 	= partial_clause_prev[493] & ~x[33] & ~x[57];
			partial_clause[494] 	= partial_clause_prev[494] & ~x[4] & ~x[27] & ~x[28] & x[50];
			partial_clause[495] 	= partial_clause_prev[495] & ~x[4] & ~x[6];
			partial_clause[496] 	= partial_clause_prev[496] & ~x[45];
			partial_clause[497] 	= partial_clause_prev[497] & 1'b1;
			partial_clause[498] 	= partial_clause_prev[498] & 1'b1;
			partial_clause[499] 	= partial_clause_prev[499] & ~x[22] & ~x[49];
		end
	end
endmodule


module HCB_4 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[52] & ~x[53];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[19] & ~x[21] & ~x[26] & ~x[46] & ~x[51];
			partial_clause[2] 	= partial_clause_prev[2] & ~x[33] & ~x[54] & ~x[57] & ~x[59];
			partial_clause[3] 	= partial_clause_prev[3] & ~x[1] & ~x[24] & ~x[37] & ~x[54];
			partial_clause[4] 	= partial_clause_prev[4] & ~x[0] & ~x[52];
			partial_clause[5] 	= partial_clause_prev[5] & ~x[20] & ~x[22] & ~x[24] & ~x[25] & ~x[29] & ~x[55] & ~x[56];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[6] & ~x[21] & ~x[32] & ~x[48] & ~x[55];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[0] & ~x[27] & ~x[28];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[1] & ~x[23] & ~x[24] & ~x[51] & ~x[53];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[23] & ~x[25] & ~x[29] & ~x[49];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[28] & ~x[49] & ~x[55];
			partial_clause[11] 	= partial_clause_prev[11] & ~x[0] & ~x[23] & ~x[26] & ~x[29] & ~x[53] & ~x[56];
			partial_clause[12] 	= partial_clause_prev[12] & ~x[1] & x[41] & ~x[47] & ~x[53] & ~x[56];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[3] & ~x[24] & ~x[25] & ~x[26] & ~x[28] & ~x[31] & ~x[58];
			partial_clause[14] 	= partial_clause_prev[14] & ~x[58];
			partial_clause[15] 	= partial_clause_prev[15] & ~x[12];
			partial_clause[16] 	= partial_clause_prev[16] & ~x[24];
			partial_clause[17] 	= partial_clause_prev[17] & 1'b1;
			partial_clause[18] 	= partial_clause_prev[18] & ~x[26] & ~x[48] & ~x[53];
			partial_clause[19] 	= partial_clause_prev[19] & ~x[48];
			partial_clause[20] 	= partial_clause_prev[20] & 1'b1;
			partial_clause[21] 	= partial_clause_prev[21] & ~x[51] & ~x[52];
			partial_clause[22] 	= partial_clause_prev[22] & ~x[25] & ~x[39] & ~x[48];
			partial_clause[23] 	= partial_clause_prev[23] & ~x[0] & ~x[7] & ~x[22] & ~x[23] & ~x[25] & ~x[26] & ~x[27] & ~x[49] & ~x[54] & ~x[55];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[0] & ~x[2] & ~x[21] & ~x[23] & ~x[25] & ~x[27] & ~x[29] & ~x[30] & ~x[50] & ~x[52] & ~x[53] & ~x[55] & ~x[57];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[0] & ~x[18] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[33] & ~x[46] & ~x[47] & ~x[49] & ~x[53] & ~x[57];
			partial_clause[26] 	= partial_clause_prev[26] & 1'b1;
			partial_clause[27] 	= partial_clause_prev[27] & ~x[2] & ~x[23] & ~x[55] & ~x[56];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[5];
			partial_clause[29] 	= partial_clause_prev[29] & ~x[23];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[50] & ~x[53] & ~x[57];
			partial_clause[31] 	= partial_clause_prev[31] & ~x[11] & ~x[13];
			partial_clause[32] 	= partial_clause_prev[32] & ~x[0] & x[37] & ~x[53] & ~x[55];
			partial_clause[33] 	= partial_clause_prev[33] & x[10];
			partial_clause[34] 	= partial_clause_prev[34] & ~x[0] & x[13] & ~x[18] & ~x[23] & ~x[24] & ~x[54] & ~x[56];
			partial_clause[35] 	= partial_clause_prev[35] & ~x[26];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[20] & ~x[50] & ~x[53];
			partial_clause[37] 	= partial_clause_prev[37] & 1'b1;
			partial_clause[38] 	= partial_clause_prev[38] & ~x[1] & ~x[3] & ~x[23] & ~x[26] & ~x[43] & ~x[44] & ~x[46] & ~x[47] & ~x[53] & ~x[60];
			partial_clause[39] 	= partial_clause_prev[39] & ~x[21] & ~x[47] & ~x[59];
			partial_clause[40] 	= partial_clause_prev[40] & ~x[21] & ~x[22] & ~x[23] & ~x[48];
			partial_clause[41] 	= partial_clause_prev[41] & 1'b1;
			partial_clause[42] 	= partial_clause_prev[42] & 1'b1;
			partial_clause[43] 	= partial_clause_prev[43] & 1'b1;
			partial_clause[44] 	= partial_clause_prev[44] & 1'b1;
			partial_clause[45] 	= partial_clause_prev[45] & ~x[24] & x[40] & ~x[45];
			partial_clause[46] 	= partial_clause_prev[46] & ~x[18] & ~x[33] & ~x[47] & ~x[48] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[54] & ~x[55] & ~x[57];
			partial_clause[47] 	= partial_clause_prev[47] & 1'b1;
			partial_clause[48] 	= partial_clause_prev[48] & 1'b1;
			partial_clause[49] 	= partial_clause_prev[49] & 1'b1;
			partial_clause[50] 	= partial_clause_prev[50] & ~x[54];
			partial_clause[51] 	= partial_clause_prev[51] & 1'b1;
			partial_clause[52] 	= partial_clause_prev[52] & 1'b1;
			partial_clause[53] 	= partial_clause_prev[53] & ~x[1] & ~x[55];
			partial_clause[54] 	= partial_clause_prev[54] & ~x[49] & ~x[52];
			partial_clause[55] 	= partial_clause_prev[55] & ~x[60];
			partial_clause[56] 	= partial_clause_prev[56] & ~x[11] & ~x[38];
			partial_clause[57] 	= partial_clause_prev[57] & x[12] & ~x[22] & ~x[26] & x[39] & ~x[45] & ~x[48];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[27] & ~x[53];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[26] & x[33] & ~x[50];
			partial_clause[60] 	= partial_clause_prev[60] & ~x[44] & ~x[50];
			partial_clause[61] 	= partial_clause_prev[61] & 1'b1;
			partial_clause[62] 	= partial_clause_prev[62] & ~x[4] & ~x[25];
			partial_clause[63] 	= partial_clause_prev[63] & ~x[17] & ~x[24] & ~x[42] & ~x[43];
			partial_clause[64] 	= partial_clause_prev[64] & 1'b1;
			partial_clause[65] 	= partial_clause_prev[65] & 1'b1;
			partial_clause[66] 	= partial_clause_prev[66] & 1'b1;
			partial_clause[67] 	= partial_clause_prev[67] & ~x[9] & ~x[35] & x[41] & ~x[61];
			partial_clause[68] 	= partial_clause_prev[68] & ~x[58];
			partial_clause[69] 	= partial_clause_prev[69] & ~x[0] & ~x[24] & ~x[51];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[28] & ~x[31] & ~x[60] & ~x[61];
			partial_clause[71] 	= partial_clause_prev[71] & ~x[21] & ~x[24];
			partial_clause[72] 	= partial_clause_prev[72] & ~x[48];
			partial_clause[73] 	= partial_clause_prev[73] & ~x[8] & ~x[36];
			partial_clause[74] 	= partial_clause_prev[74] & ~x[23] & ~x[46] & ~x[50];
			partial_clause[75] 	= partial_clause_prev[75] & 1'b1;
			partial_clause[76] 	= partial_clause_prev[76] & ~x[12] & ~x[24] & ~x[29] & ~x[49] & ~x[58];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[3] & ~x[14] & ~x[16] & ~x[17] & ~x[41] & ~x[49];
			partial_clause[78] 	= partial_clause_prev[78] & ~x[60];
			partial_clause[79] 	= partial_clause_prev[79] & ~x[28] & ~x[47] & ~x[51];
			partial_clause[80] 	= partial_clause_prev[80] & ~x[39];
			partial_clause[81] 	= partial_clause_prev[81] & 1'b1;
			partial_clause[82] 	= partial_clause_prev[82] & ~x[3] & ~x[23];
			partial_clause[83] 	= partial_clause_prev[83] & ~x[59];
			partial_clause[84] 	= partial_clause_prev[84] & x[10] & ~x[55];
			partial_clause[85] 	= partial_clause_prev[85] & ~x[1] & ~x[53] & ~x[57];
			partial_clause[86] 	= partial_clause_prev[86] & ~x[21] & ~x[28] & ~x[55];
			partial_clause[87] 	= partial_clause_prev[87] & ~x[12] & ~x[14] & ~x[15] & ~x[23] & ~x[43] & ~x[49];
			partial_clause[88] 	= partial_clause_prev[88] & ~x[23] & ~x[27] & ~x[50] & ~x[52] & ~x[53];
			partial_clause[89] 	= partial_clause_prev[89] & x[10] & x[11];
			partial_clause[90] 	= partial_clause_prev[90] & ~x[11];
			partial_clause[91] 	= partial_clause_prev[91] & x[14];
			partial_clause[92] 	= partial_clause_prev[92] & ~x[44] & ~x[45] & ~x[54];
			partial_clause[93] 	= partial_clause_prev[93] & ~x[17] & ~x[22] & ~x[26] & ~x[27] & ~x[38] & ~x[47] & ~x[49] & ~x[51] & ~x[54] & ~x[55] & ~x[56];
			partial_clause[94] 	= partial_clause_prev[94] & x[9];
			partial_clause[95] 	= partial_clause_prev[95] & ~x[1] & ~x[2] & ~x[20] & ~x[31] & ~x[49];
			partial_clause[96] 	= partial_clause_prev[96] & 1'b1;
			partial_clause[97] 	= partial_clause_prev[97] & ~x[0] & ~x[1] & ~x[19] & ~x[23] & ~x[25] & ~x[26] & ~x[28] & ~x[49] & ~x[54];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[0] & ~x[1] & ~x[2] & ~x[24] & ~x[27] & ~x[28] & ~x[29] & ~x[46] & ~x[52] & ~x[54] & ~x[56];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[0] & ~x[20] & ~x[25] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[55];
			partial_clause[100] 	= partial_clause_prev[100] & ~x[2] & ~x[19] & ~x[48];
			partial_clause[101] 	= partial_clause_prev[101] & 1'b1;
			partial_clause[102] 	= partial_clause_prev[102] & ~x[4] & ~x[51] & ~x[53];
			partial_clause[103] 	= partial_clause_prev[103] & ~x[18] & ~x[22] & ~x[23] & ~x[27] & ~x[28] & ~x[29] & ~x[46] & ~x[48] & ~x[49] & ~x[50] & ~x[52] & ~x[57];
			partial_clause[104] 	= partial_clause_prev[104] & ~x[22] & ~x[29];
			partial_clause[105] 	= partial_clause_prev[105] & ~x[20] & ~x[22] & ~x[50] & ~x[53];
			partial_clause[106] 	= partial_clause_prev[106] & ~x[27] & ~x[54];
			partial_clause[107] 	= partial_clause_prev[107] & ~x[0] & ~x[21] & ~x[22] & ~x[28] & ~x[29] & ~x[52] & ~x[56];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[49];
			partial_clause[109] 	= partial_clause_prev[109] & ~x[10] & ~x[37];
			partial_clause[110] 	= partial_clause_prev[110] & 1'b1;
			partial_clause[111] 	= partial_clause_prev[111] & x[60];
			partial_clause[112] 	= partial_clause_prev[112] & ~x[14] & ~x[15] & ~x[20];
			partial_clause[113] 	= partial_clause_prev[113] & ~x[20];
			partial_clause[114] 	= partial_clause_prev[114] & 1'b1;
			partial_clause[115] 	= partial_clause_prev[115] & ~x[49] & ~x[52] & ~x[53] & ~x[55];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[1] & ~x[51] & ~x[56];
			partial_clause[117] 	= partial_clause_prev[117] & ~x[6] & ~x[31] & ~x[59];
			partial_clause[118] 	= partial_clause_prev[118] & 1'b1;
			partial_clause[119] 	= partial_clause_prev[119] & ~x[26] & ~x[47] & ~x[48] & ~x[53];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[0] & ~x[21] & ~x[23] & ~x[28] & ~x[52] & ~x[54] & ~x[56];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[28] & ~x[52];
			partial_clause[122] 	= partial_clause_prev[122] & ~x[31] & ~x[53] & ~x[55];
			partial_clause[123] 	= partial_clause_prev[123] & ~x[0] & ~x[1] & ~x[2] & ~x[4] & ~x[21] & ~x[28] & ~x[33] & ~x[42] & ~x[45] & ~x[47] & ~x[48] & ~x[49] & ~x[58] & ~x[60];
			partial_clause[124] 	= partial_clause_prev[124] & ~x[55];
			partial_clause[125] 	= partial_clause_prev[125] & ~x[30];
			partial_clause[126] 	= partial_clause_prev[126] & 1'b1;
			partial_clause[127] 	= partial_clause_prev[127] & ~x[0] & ~x[51] & ~x[52] & ~x[53] & ~x[54] & ~x[55];
			partial_clause[128] 	= partial_clause_prev[128] & x[6];
			partial_clause[129] 	= partial_clause_prev[129] & ~x[4] & ~x[21] & ~x[24] & ~x[27] & ~x[29] & ~x[32] & x[36] & ~x[48] & ~x[49] & ~x[51] & ~x[52] & ~x[55];
			partial_clause[130] 	= partial_clause_prev[130] & ~x[19] & ~x[20] & ~x[22] & ~x[25] & ~x[28] & ~x[47] & ~x[50] & ~x[52] & ~x[54];
			partial_clause[131] 	= partial_clause_prev[131] & x[41] & ~x[53];
			partial_clause[132] 	= partial_clause_prev[132] & ~x[3] & ~x[4] & ~x[16] & ~x[30] & ~x[44] & ~x[49] & ~x[52] & ~x[60];
			partial_clause[133] 	= partial_clause_prev[133] & ~x[22];
			partial_clause[134] 	= partial_clause_prev[134] & ~x[23] & ~x[26] & ~x[28] & ~x[49] & ~x[50] & ~x[53] & ~x[54];
			partial_clause[135] 	= partial_clause_prev[135] & ~x[2];
			partial_clause[136] 	= partial_clause_prev[136] & ~x[22] & ~x[27] & ~x[28] & ~x[51];
			partial_clause[137] 	= partial_clause_prev[137] & ~x[21];
			partial_clause[138] 	= partial_clause_prev[138] & 1'b1;
			partial_clause[139] 	= partial_clause_prev[139] & ~x[18] & ~x[47] & ~x[53] & ~x[56] & ~x[59];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[2] & ~x[4] & ~x[19] & ~x[25] & ~x[48] & ~x[50] & ~x[51] & ~x[54] & ~x[56] & ~x[59];
			partial_clause[141] 	= partial_clause_prev[141] & ~x[16] & ~x[21];
			partial_clause[142] 	= partial_clause_prev[142] & ~x[0] & ~x[1] & ~x[25] & ~x[27] & ~x[28] & ~x[38] & ~x[52] & ~x[54];
			partial_clause[143] 	= partial_clause_prev[143] & ~x[53];
			partial_clause[144] 	= partial_clause_prev[144] & ~x[0] & ~x[53];
			partial_clause[145] 	= partial_clause_prev[145] & ~x[28] & x[34];
			partial_clause[146] 	= partial_clause_prev[146] & ~x[54] & ~x[55];
			partial_clause[147] 	= partial_clause_prev[147] & ~x[0] & ~x[30] & ~x[44] & ~x[48] & ~x[51] & ~x[53] & ~x[56];
			partial_clause[148] 	= partial_clause_prev[148] & ~x[22];
			partial_clause[149] 	= partial_clause_prev[149] & ~x[2] & ~x[51];
			partial_clause[150] 	= partial_clause_prev[150] & ~x[21] & ~x[24] & ~x[26] & ~x[28] & ~x[31] & ~x[53];
			partial_clause[151] 	= partial_clause_prev[151] & 1'b1;
			partial_clause[152] 	= partial_clause_prev[152] & ~x[27];
			partial_clause[153] 	= partial_clause_prev[153] & ~x[20] & ~x[27] & ~x[48] & ~x[51] & ~x[55];
			partial_clause[154] 	= partial_clause_prev[154] & ~x[56];
			partial_clause[155] 	= partial_clause_prev[155] & 1'b1;
			partial_clause[156] 	= partial_clause_prev[156] & 1'b1;
			partial_clause[157] 	= partial_clause_prev[157] & 1'b1;
			partial_clause[158] 	= partial_clause_prev[158] & ~x[22] & ~x[23] & ~x[25] & ~x[27] & ~x[29] & ~x[50] & ~x[51] & ~x[53] & ~x[54] & ~x[55] & ~x[56];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[25] & ~x[32] & ~x[48] & ~x[51] & ~x[55];
			partial_clause[160] 	= partial_clause_prev[160] & ~x[43] & ~x[44] & ~x[52];
			partial_clause[161] 	= partial_clause_prev[161] & ~x[24] & ~x[34] & ~x[49] & ~x[57] & ~x[60];
			partial_clause[162] 	= partial_clause_prev[162] & ~x[23] & ~x[50];
			partial_clause[163] 	= partial_clause_prev[163] & x[38];
			partial_clause[164] 	= partial_clause_prev[164] & ~x[22] & ~x[27];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[26] & ~x[47] & ~x[50] & ~x[52];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[26] & ~x[54] & ~x[55];
			partial_clause[167] 	= partial_clause_prev[167] & ~x[11] & ~x[39];
			partial_clause[168] 	= partial_clause_prev[168] & 1'b1;
			partial_clause[169] 	= partial_clause_prev[169] & 1'b1;
			partial_clause[170] 	= partial_clause_prev[170] & ~x[21];
			partial_clause[171] 	= partial_clause_prev[171] & ~x[22] & ~x[51];
			partial_clause[172] 	= partial_clause_prev[172] & x[12];
			partial_clause[173] 	= partial_clause_prev[173] & x[16] & ~x[20] & ~x[21];
			partial_clause[174] 	= partial_clause_prev[174] & ~x[24];
			partial_clause[175] 	= partial_clause_prev[175] & ~x[57] & ~x[59];
			partial_clause[176] 	= partial_clause_prev[176] & ~x[59] & ~x[62];
			partial_clause[177] 	= partial_clause_prev[177] & ~x[20];
			partial_clause[178] 	= partial_clause_prev[178] & ~x[24] & ~x[38];
			partial_clause[179] 	= partial_clause_prev[179] & ~x[11] & ~x[39];
			partial_clause[180] 	= partial_clause_prev[180] & ~x[56];
			partial_clause[181] 	= partial_clause_prev[181] & 1'b1;
			partial_clause[182] 	= partial_clause_prev[182] & 1'b1;
			partial_clause[183] 	= partial_clause_prev[183] & ~x[0] & ~x[2] & ~x[26] & ~x[30] & ~x[57];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[27] & ~x[30] & ~x[31] & ~x[51] & ~x[52] & ~x[56];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[1] & ~x[29];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[2] & ~x[31] & ~x[46] & ~x[50];
			partial_clause[187] 	= partial_clause_prev[187] & ~x[19] & ~x[25] & ~x[49] & ~x[54];
			partial_clause[188] 	= partial_clause_prev[188] & ~x[50] & ~x[55];
			partial_clause[189] 	= partial_clause_prev[189] & 1'b1;
			partial_clause[190] 	= partial_clause_prev[190] & ~x[1] & ~x[24] & ~x[55];
			partial_clause[191] 	= partial_clause_prev[191] & ~x[6] & ~x[17] & ~x[21] & ~x[47] & ~x[48] & ~x[51] & ~x[57] & ~x[59];
			partial_clause[192] 	= partial_clause_prev[192] & ~x[41] & ~x[44] & ~x[45] & ~x[47];
			partial_clause[193] 	= partial_clause_prev[193] & ~x[16] & ~x[18] & ~x[25] & ~x[29];
			partial_clause[194] 	= partial_clause_prev[194] & ~x[42];
			partial_clause[195] 	= partial_clause_prev[195] & ~x[26] & ~x[30] & ~x[53];
			partial_clause[196] 	= partial_clause_prev[196] & ~x[47];
			partial_clause[197] 	= partial_clause_prev[197] & ~x[3] & ~x[19] & ~x[25] & ~x[47] & ~x[48] & ~x[49] & ~x[53] & ~x[56] & ~x[58] & ~x[59];
			partial_clause[198] 	= partial_clause_prev[198] & x[8] & x[13] & x[14];
			partial_clause[199] 	= partial_clause_prev[199] & 1'b1;
			partial_clause[200] 	= partial_clause_prev[200] & ~x[21] & ~x[50];
			partial_clause[201] 	= partial_clause_prev[201] & ~x[6] & ~x[27] & ~x[60];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[0] & ~x[19] & ~x[29] & ~x[49] & ~x[56];
			partial_clause[203] 	= partial_clause_prev[203] & 1'b1;
			partial_clause[204] 	= partial_clause_prev[204] & ~x[0] & ~x[3] & ~x[4] & ~x[24] & ~x[25] & ~x[26] & ~x[49] & ~x[50] & ~x[51] & ~x[52] & ~x[54];
			partial_clause[205] 	= partial_clause_prev[205] & ~x[26];
			partial_clause[206] 	= partial_clause_prev[206] & 1'b1;
			partial_clause[207] 	= partial_clause_prev[207] & ~x[1] & ~x[17] & ~x[26] & ~x[44] & ~x[45] & ~x[56] & ~x[57];
			partial_clause[208] 	= partial_clause_prev[208] & x[41] & ~x[53] & ~x[54];
			partial_clause[209] 	= partial_clause_prev[209] & ~x[33] & ~x[58];
			partial_clause[210] 	= partial_clause_prev[210] & ~x[4] & ~x[6] & ~x[7] & ~x[8] & ~x[21] & ~x[24] & ~x[30] & ~x[48] & ~x[49] & ~x[56] & ~x[58];
			partial_clause[211] 	= partial_clause_prev[211] & ~x[2] & ~x[7];
			partial_clause[212] 	= partial_clause_prev[212] & ~x[17] & ~x[29] & ~x[49];
			partial_clause[213] 	= partial_clause_prev[213] & 1'b1;
			partial_clause[214] 	= partial_clause_prev[214] & ~x[0];
			partial_clause[215] 	= partial_clause_prev[215] & ~x[0] & ~x[3] & ~x[18] & ~x[31] & ~x[48];
			partial_clause[216] 	= partial_clause_prev[216] & ~x[49];
			partial_clause[217] 	= partial_clause_prev[217] & ~x[11] & ~x[19] & ~x[20] & ~x[26] & ~x[49] & ~x[50] & ~x[51];
			partial_clause[218] 	= partial_clause_prev[218] & x[11] & ~x[28];
			partial_clause[219] 	= partial_clause_prev[219] & ~x[19] & ~x[20] & ~x[47];
			partial_clause[220] 	= partial_clause_prev[220] & ~x[25] & ~x[53] & ~x[55];
			partial_clause[221] 	= partial_clause_prev[221] & ~x[47];
			partial_clause[222] 	= partial_clause_prev[222] & ~x[4] & x[63];
			partial_clause[223] 	= partial_clause_prev[223] & ~x[29] & ~x[51] & ~x[53];
			partial_clause[224] 	= partial_clause_prev[224] & ~x[3] & ~x[21] & ~x[28] & ~x[29] & ~x[30] & ~x[49] & ~x[56] & ~x[58];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[21] & ~x[22] & ~x[23] & ~x[53] & ~x[54] & ~x[55];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[23] & ~x[25] & ~x[26] & ~x[28] & ~x[50] & ~x[51];
			partial_clause[227] 	= partial_clause_prev[227] & ~x[19] & ~x[20] & ~x[26] & ~x[49] & ~x[51] & ~x[53] & ~x[54];
			partial_clause[228] 	= partial_clause_prev[228] & ~x[1] & ~x[22] & ~x[32] & x[35] & ~x[51] & ~x[53] & ~x[54] & ~x[58] & ~x[60];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[1] & ~x[3] & ~x[52] & ~x[53] & ~x[56];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[1] & ~x[25] & ~x[26] & ~x[27] & ~x[52];
			partial_clause[231] 	= partial_clause_prev[231] & ~x[1] & ~x[22] & ~x[50];
			partial_clause[232] 	= partial_clause_prev[232] & 1'b1;
			partial_clause[233] 	= partial_clause_prev[233] & ~x[52] & ~x[62];
			partial_clause[234] 	= partial_clause_prev[234] & ~x[50];
			partial_clause[235] 	= partial_clause_prev[235] & 1'b1;
			partial_clause[236] 	= partial_clause_prev[236] & 1'b1;
			partial_clause[237] 	= partial_clause_prev[237] & ~x[34];
			partial_clause[238] 	= partial_clause_prev[238] & ~x[53];
			partial_clause[239] 	= partial_clause_prev[239] & ~x[28];
			partial_clause[240] 	= partial_clause_prev[240] & ~x[31] & ~x[51] & ~x[59];
			partial_clause[241] 	= partial_clause_prev[241] & ~x[49];
			partial_clause[242] 	= partial_clause_prev[242] & ~x[26] & ~x[54] & ~x[56] & ~x[58];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[20] & ~x[22] & ~x[24] & ~x[36] & ~x[37] & ~x[50] & ~x[52] & ~x[53] & ~x[55];
			partial_clause[244] 	= partial_clause_prev[244] & ~x[10] & ~x[22] & ~x[26];
			partial_clause[245] 	= partial_clause_prev[245] & 1'b1;
			partial_clause[246] 	= partial_clause_prev[246] & ~x[26];
			partial_clause[247] 	= partial_clause_prev[247] & ~x[26] & ~x[27] & ~x[39] & ~x[49] & ~x[50] & ~x[53];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[0] & ~x[1] & ~x[9] & ~x[17] & ~x[21] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & ~x[48] & ~x[51] & ~x[52] & ~x[53] & ~x[55] & ~x[56];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[18] & ~x[19] & ~x[44] & ~x[47];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[0] & ~x[23] & ~x[25] & ~x[26] & ~x[27] & ~x[29] & ~x[50] & ~x[51] & ~x[53] & ~x[54] & ~x[55] & ~x[58];
			partial_clause[251] 	= partial_clause_prev[251] & ~x[3] & ~x[26];
			partial_clause[252] 	= partial_clause_prev[252] & ~x[0] & ~x[9] & ~x[22] & ~x[50] & ~x[52] & ~x[53];
			partial_clause[253] 	= partial_clause_prev[253] & x[10] & ~x[23] & ~x[26];
			partial_clause[254] 	= partial_clause_prev[254] & ~x[0] & ~x[10] & ~x[18] & ~x[24] & ~x[51];
			partial_clause[255] 	= partial_clause_prev[255] & ~x[24] & ~x[47] & ~x[56];
			partial_clause[256] 	= partial_clause_prev[256] & 1'b1;
			partial_clause[257] 	= partial_clause_prev[257] & ~x[22] & ~x[53];
			partial_clause[258] 	= partial_clause_prev[258] & ~x[51] & ~x[52];
			partial_clause[259] 	= partial_clause_prev[259] & 1'b1;
			partial_clause[260] 	= partial_clause_prev[260] & ~x[50];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[21] & ~x[24] & ~x[26] & ~x[29] & ~x[52] & ~x[57];
			partial_clause[262] 	= partial_clause_prev[262] & ~x[1] & ~x[47];
			partial_clause[263] 	= partial_clause_prev[263] & ~x[22];
			partial_clause[264] 	= partial_clause_prev[264] & ~x[4];
			partial_clause[265] 	= partial_clause_prev[265] & 1'b1;
			partial_clause[266] 	= partial_clause_prev[266] & ~x[21] & ~x[23];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[24] & ~x[25] & ~x[50] & ~x[52] & ~x[55];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[0] & ~x[21] & ~x[28] & ~x[51] & ~x[56] & ~x[58];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[0] & ~x[1] & ~x[24] & ~x[25] & ~x[40] & ~x[52] & ~x[53] & ~x[56];
			partial_clause[270] 	= partial_clause_prev[270] & x[38];
			partial_clause[271] 	= partial_clause_prev[271] & ~x[50] & ~x[55];
			partial_clause[272] 	= partial_clause_prev[272] & ~x[39] & ~x[48];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[27] & ~x[49] & ~x[51] & ~x[53] & ~x[55];
			partial_clause[274] 	= partial_clause_prev[274] & ~x[7] & ~x[21] & ~x[33] & ~x[34];
			partial_clause[275] 	= partial_clause_prev[275] & 1'b1;
			partial_clause[276] 	= partial_clause_prev[276] & ~x[24] & ~x[50] & ~x[56];
			partial_clause[277] 	= partial_clause_prev[277] & ~x[41] & ~x[51] & ~x[53];
			partial_clause[278] 	= partial_clause_prev[278] & 1'b1;
			partial_clause[279] 	= partial_clause_prev[279] & ~x[1] & ~x[26] & ~x[47] & ~x[55];
			partial_clause[280] 	= partial_clause_prev[280] & 1'b1;
			partial_clause[281] 	= partial_clause_prev[281] & ~x[14] & ~x[20] & ~x[26] & ~x[27] & ~x[49] & ~x[55] & ~x[59];
			partial_clause[282] 	= partial_clause_prev[282] & ~x[30];
			partial_clause[283] 	= partial_clause_prev[283] & ~x[24] & ~x[48] & ~x[52];
			partial_clause[284] 	= partial_clause_prev[284] & ~x[60];
			partial_clause[285] 	= partial_clause_prev[285] & 1'b1;
			partial_clause[286] 	= partial_clause_prev[286] & ~x[26];
			partial_clause[287] 	= partial_clause_prev[287] & ~x[24] & ~x[51];
			partial_clause[288] 	= partial_clause_prev[288] & 1'b1;
			partial_clause[289] 	= partial_clause_prev[289] & ~x[7] & ~x[34];
			partial_clause[290] 	= partial_clause_prev[290] & ~x[8] & ~x[9] & ~x[55] & ~x[59];
			partial_clause[291] 	= partial_clause_prev[291] & x[12] & ~x[30];
			partial_clause[292] 	= partial_clause_prev[292] & ~x[26] & ~x[48];
			partial_clause[293] 	= partial_clause_prev[293] & ~x[50];
			partial_clause[294] 	= partial_clause_prev[294] & 1'b1;
			partial_clause[295] 	= partial_clause_prev[295] & 1'b1;
			partial_clause[296] 	= partial_clause_prev[296] & x[41] & ~x[56] & ~x[58];
			partial_clause[297] 	= partial_clause_prev[297] & ~x[24] & ~x[27];
			partial_clause[298] 	= partial_clause_prev[298] & ~x[11] & ~x[12] & ~x[14] & ~x[18] & ~x[43] & ~x[44] & ~x[45];
			partial_clause[299] 	= partial_clause_prev[299] & ~x[5] & ~x[19] & ~x[33] & x[37] & ~x[46] & ~x[55];
			partial_clause[300] 	= partial_clause_prev[300] & ~x[21];
			partial_clause[301] 	= partial_clause_prev[301] & ~x[1] & ~x[20] & ~x[24] & ~x[29];
			partial_clause[302] 	= partial_clause_prev[302] & 1'b1;
			partial_clause[303] 	= partial_clause_prev[303] & 1'b1;
			partial_clause[304] 	= partial_clause_prev[304] & ~x[10] & ~x[31] & ~x[36] & ~x[58] & ~x[61];
			partial_clause[305] 	= partial_clause_prev[305] & 1'b1;
			partial_clause[306] 	= partial_clause_prev[306] & ~x[1] & ~x[22] & ~x[40] & ~x[52] & ~x[54] & ~x[55];
			partial_clause[307] 	= partial_clause_prev[307] & ~x[19] & ~x[28] & ~x[46] & ~x[47] & ~x[57];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[17] & ~x[46];
			partial_clause[309] 	= partial_clause_prev[309] & 1'b1;
			partial_clause[310] 	= partial_clause_prev[310] & 1'b1;
			partial_clause[311] 	= partial_clause_prev[311] & ~x[24] & ~x[26];
			partial_clause[312] 	= partial_clause_prev[312] & ~x[22] & ~x[52];
			partial_clause[313] 	= partial_clause_prev[313] & ~x[49];
			partial_clause[314] 	= partial_clause_prev[314] & 1'b1;
			partial_clause[315] 	= partial_clause_prev[315] & ~x[24] & ~x[25];
			partial_clause[316] 	= partial_clause_prev[316] & ~x[24] & ~x[27];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[19];
			partial_clause[318] 	= partial_clause_prev[318] & ~x[2] & ~x[30] & ~x[49] & ~x[60];
			partial_clause[319] 	= partial_clause_prev[319] & ~x[25] & ~x[54] & ~x[58];
			partial_clause[320] 	= partial_clause_prev[320] & ~x[0] & ~x[52];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[24] & ~x[29] & ~x[53] & ~x[54] & ~x[56];
			partial_clause[322] 	= partial_clause_prev[322] & 1'b1;
			partial_clause[323] 	= partial_clause_prev[323] & x[7] & x[9] & x[11];
			partial_clause[324] 	= partial_clause_prev[324] & ~x[26] & ~x[42];
			partial_clause[325] 	= partial_clause_prev[325] & ~x[2] & ~x[24] & ~x[26] & ~x[29] & ~x[51] & ~x[53];
			partial_clause[326] 	= partial_clause_prev[326] & ~x[25] & ~x[50] & ~x[52] & ~x[54] & ~x[56] & x[59];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[0] & ~x[24] & ~x[26] & ~x[57];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[25] & ~x[50] & ~x[55] & ~x[59];
			partial_clause[329] 	= partial_clause_prev[329] & x[42];
			partial_clause[330] 	= partial_clause_prev[330] & 1'b1;
			partial_clause[331] 	= partial_clause_prev[331] & ~x[31] & ~x[57];
			partial_clause[332] 	= partial_clause_prev[332] & ~x[0] & ~x[28] & ~x[45] & ~x[50] & ~x[55];
			partial_clause[333] 	= partial_clause_prev[333] & ~x[21] & ~x[24] & ~x[35] & ~x[37] & ~x[61];
			partial_clause[334] 	= partial_clause_prev[334] & 1'b1;
			partial_clause[335] 	= partial_clause_prev[335] & ~x[49] & ~x[63];
			partial_clause[336] 	= partial_clause_prev[336] & x[13];
			partial_clause[337] 	= partial_clause_prev[337] & ~x[3] & ~x[20] & ~x[23] & ~x[31] & ~x[56] & ~x[59];
			partial_clause[338] 	= partial_clause_prev[338] & ~x[29];
			partial_clause[339] 	= partial_clause_prev[339] & ~x[27] & ~x[28] & ~x[51];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[19] & ~x[22] & ~x[23];
			partial_clause[341] 	= partial_clause_prev[341] & ~x[34] & ~x[36];
			partial_clause[342] 	= partial_clause_prev[342] & ~x[49] & ~x[54];
			partial_clause[343] 	= partial_clause_prev[343] & x[12] & ~x[19] & ~x[22] & ~x[23] & ~x[26] & ~x[48] & ~x[52];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[16] & ~x[22] & ~x[31] & ~x[44];
			partial_clause[345] 	= partial_clause_prev[345] & ~x[5] & ~x[6] & ~x[30];
			partial_clause[346] 	= partial_clause_prev[346] & ~x[49] & ~x[51] & ~x[52];
			partial_clause[347] 	= partial_clause_prev[347] & ~x[22] & ~x[25] & ~x[50] & ~x[51] & ~x[55];
			partial_clause[348] 	= partial_clause_prev[348] & ~x[20] & ~x[54];
			partial_clause[349] 	= partial_clause_prev[349] & ~x[55];
			partial_clause[350] 	= partial_clause_prev[350] & ~x[0] & ~x[17] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[25] & ~x[26] & ~x[28] & ~x[44] & ~x[51] & ~x[52] & ~x[53] & ~x[54];
			partial_clause[351] 	= partial_clause_prev[351] & 1'b1;
			partial_clause[352] 	= partial_clause_prev[352] & 1'b1;
			partial_clause[353] 	= partial_clause_prev[353] & 1'b1;
			partial_clause[354] 	= partial_clause_prev[354] & ~x[5] & ~x[8] & ~x[22] & ~x[37] & ~x[60];
			partial_clause[355] 	= partial_clause_prev[355] & ~x[35];
			partial_clause[356] 	= partial_clause_prev[356] & ~x[0] & ~x[48];
			partial_clause[357] 	= partial_clause_prev[357] & ~x[25] & x[33];
			partial_clause[358] 	= partial_clause_prev[358] & ~x[25] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[54] & ~x[55] & ~x[56];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[9] & ~x[53] & ~x[54];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[19] & ~x[48] & ~x[49] & ~x[51] & ~x[53];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[1] & ~x[40] & ~x[56];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[51];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[2] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[25] & ~x[31] & ~x[44] & ~x[51] & ~x[58];
			partial_clause[364] 	= partial_clause_prev[364] & ~x[20] & ~x[24] & ~x[48] & ~x[58];
			partial_clause[365] 	= partial_clause_prev[365] & x[32] & ~x[35];
			partial_clause[366] 	= partial_clause_prev[366] & ~x[24] & ~x[25] & ~x[49] & ~x[50] & ~x[51] & ~x[53] & ~x[55];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[22] & ~x[41];
			partial_clause[368] 	= partial_clause_prev[368] & ~x[9] & ~x[11];
			partial_clause[369] 	= partial_clause_prev[369] & ~x[49] & ~x[52];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[18] & ~x[20] & ~x[23] & ~x[51] & ~x[53];
			partial_clause[371] 	= partial_clause_prev[371] & ~x[42] & ~x[44];
			partial_clause[372] 	= partial_clause_prev[372] & ~x[21];
			partial_clause[373] 	= partial_clause_prev[373] & 1'b1;
			partial_clause[374] 	= partial_clause_prev[374] & ~x[49];
			partial_clause[375] 	= partial_clause_prev[375] & 1'b1;
			partial_clause[376] 	= partial_clause_prev[376] & ~x[28] & ~x[47] & ~x[53] & ~x[56] & ~x[58];
			partial_clause[377] 	= partial_clause_prev[377] & ~x[20] & ~x[21] & ~x[50];
			partial_clause[378] 	= partial_clause_prev[378] & ~x[1] & ~x[13] & ~x[43] & ~x[58];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[22] & ~x[38] & ~x[62] & ~x[63];
			partial_clause[380] 	= partial_clause_prev[380] & ~x[39] & ~x[56];
			partial_clause[381] 	= partial_clause_prev[381] & ~x[10] & ~x[22] & ~x[25] & ~x[48] & ~x[54] & ~x[55];
			partial_clause[382] 	= partial_clause_prev[382] & 1'b1;
			partial_clause[383] 	= partial_clause_prev[383] & ~x[7] & ~x[34];
			partial_clause[384] 	= partial_clause_prev[384] & ~x[39] & ~x[41] & ~x[42] & ~x[45] & ~x[47];
			partial_clause[385] 	= partial_clause_prev[385] & 1'b1;
			partial_clause[386] 	= partial_clause_prev[386] & 1'b1;
			partial_clause[387] 	= partial_clause_prev[387] & ~x[29] & ~x[52] & ~x[55] & ~x[57];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[22] & ~x[24] & ~x[26] & ~x[27] & ~x[39] & ~x[53] & ~x[54];
			partial_clause[389] 	= partial_clause_prev[389] & ~x[4] & ~x[40];
			partial_clause[390] 	= partial_clause_prev[390] & ~x[9] & ~x[20] & ~x[21] & ~x[26] & ~x[47] & ~x[53];
			partial_clause[391] 	= partial_clause_prev[391] & ~x[9];
			partial_clause[392] 	= partial_clause_prev[392] & ~x[48];
			partial_clause[393] 	= partial_clause_prev[393] & ~x[6] & ~x[8] & ~x[31];
			partial_clause[394] 	= partial_clause_prev[394] & ~x[18] & ~x[25] & ~x[31] & ~x[34] & ~x[36] & ~x[47] & ~x[60];
			partial_clause[395] 	= partial_clause_prev[395] & ~x[0] & x[35] & ~x[55] & x[63];
			partial_clause[396] 	= partial_clause_prev[396] & ~x[57];
			partial_clause[397] 	= partial_clause_prev[397] & 1'b1;
			partial_clause[398] 	= partial_clause_prev[398] & ~x[40] & ~x[41];
			partial_clause[399] 	= partial_clause_prev[399] & 1'b1;
			partial_clause[400] 	= partial_clause_prev[400] & ~x[19] & ~x[20] & ~x[23] & ~x[49];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[24] & ~x[26] & ~x[27] & ~x[30] & ~x[50];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[20] & ~x[48] & ~x[51] & ~x[53] & ~x[54];
			partial_clause[403] 	= partial_clause_prev[403] & ~x[52];
			partial_clause[404] 	= partial_clause_prev[404] & 1'b1;
			partial_clause[405] 	= partial_clause_prev[405] & ~x[1];
			partial_clause[406] 	= partial_clause_prev[406] & ~x[24] & ~x[49];
			partial_clause[407] 	= partial_clause_prev[407] & x[36];
			partial_clause[408] 	= partial_clause_prev[408] & ~x[21] & ~x[27] & ~x[28] & x[33];
			partial_clause[409] 	= partial_clause_prev[409] & ~x[1] & ~x[18] & ~x[21] & ~x[22] & ~x[23] & ~x[26] & ~x[29] & ~x[46] & ~x[48] & ~x[50] & ~x[54];
			partial_clause[410] 	= partial_clause_prev[410] & ~x[44] & ~x[48];
			partial_clause[411] 	= partial_clause_prev[411] & ~x[0] & ~x[3] & ~x[19] & ~x[46] & ~x[50] & ~x[51] & ~x[53];
			partial_clause[412] 	= partial_clause_prev[412] & ~x[1] & ~x[3] & ~x[22] & ~x[23] & ~x[26] & ~x[31] & ~x[32] & ~x[49] & ~x[53] & ~x[54] & ~x[55];
			partial_clause[413] 	= partial_clause_prev[413] & ~x[1] & ~x[20] & ~x[22] & ~x[24] & ~x[49] & ~x[52];
			partial_clause[414] 	= partial_clause_prev[414] & ~x[0] & ~x[2] & ~x[29] & ~x[53] & ~x[56];
			partial_clause[415] 	= partial_clause_prev[415] & ~x[7] & ~x[16] & ~x[19] & ~x[20] & ~x[33] & ~x[46] & ~x[54] & ~x[55] & ~x[57] & ~x[59];
			partial_clause[416] 	= partial_clause_prev[416] & ~x[22] & ~x[28] & ~x[54] & ~x[55];
			partial_clause[417] 	= partial_clause_prev[417] & ~x[20] & ~x[32] & ~x[52];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[1] & ~x[2] & ~x[24] & ~x[26] & ~x[28] & ~x[30] & ~x[47] & ~x[52] & ~x[54] & ~x[56] & ~x[57];
			partial_clause[419] 	= partial_clause_prev[419] & ~x[20] & ~x[31] & ~x[37] & ~x[61] & ~x[63];
			partial_clause[420] 	= partial_clause_prev[420] & 1'b1;
			partial_clause[421] 	= partial_clause_prev[421] & ~x[25];
			partial_clause[422] 	= partial_clause_prev[422] & ~x[53];
			partial_clause[423] 	= partial_clause_prev[423] & ~x[28];
			partial_clause[424] 	= partial_clause_prev[424] & ~x[5] & ~x[50];
			partial_clause[425] 	= partial_clause_prev[425] & ~x[57];
			partial_clause[426] 	= partial_clause_prev[426] & ~x[23] & ~x[24] & ~x[29] & ~x[50] & ~x[56] & ~x[57];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[22] & ~x[23] & ~x[24] & ~x[56];
			partial_clause[428] 	= partial_clause_prev[428] & 1'b1;
			partial_clause[429] 	= partial_clause_prev[429] & 1'b1;
			partial_clause[430] 	= partial_clause_prev[430] & ~x[0] & ~x[3] & ~x[22] & ~x[50] & ~x[55] & ~x[62];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[31] & ~x[33] & ~x[47] & ~x[58] & ~x[59];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[50] & ~x[51] & ~x[52];
			partial_clause[433] 	= partial_clause_prev[433] & ~x[51] & ~x[54];
			partial_clause[434] 	= partial_clause_prev[434] & 1'b1;
			partial_clause[435] 	= partial_clause_prev[435] & ~x[0] & ~x[19] & ~x[20] & ~x[27] & ~x[28] & ~x[49] & ~x[54] & ~x[55];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[8] & ~x[9] & ~x[19] & ~x[21] & ~x[25] & ~x[35] & ~x[58] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[3] & ~x[4] & x[8] & ~x[32] & ~x[55] & ~x[56];
			partial_clause[438] 	= partial_clause_prev[438] & ~x[26];
			partial_clause[439] 	= partial_clause_prev[439] & ~x[3] & ~x[9] & ~x[28] & ~x[35] & ~x[47] & ~x[48] & ~x[51] & ~x[55] & ~x[56] & ~x[61];
			partial_clause[440] 	= partial_clause_prev[440] & ~x[29];
			partial_clause[441] 	= partial_clause_prev[441] & ~x[0] & ~x[11] & ~x[26] & ~x[51] & ~x[53] & ~x[54];
			partial_clause[442] 	= partial_clause_prev[442] & 1'b1;
			partial_clause[443] 	= partial_clause_prev[443] & ~x[0] & ~x[26] & ~x[47] & ~x[49] & ~x[57];
			partial_clause[444] 	= partial_clause_prev[444] & x[15];
			partial_clause[445] 	= partial_clause_prev[445] & 1'b1;
			partial_clause[446] 	= partial_clause_prev[446] & ~x[25] & ~x[46] & ~x[51] & ~x[52] & ~x[53];
			partial_clause[447] 	= partial_clause_prev[447] & ~x[24] & ~x[51] & ~x[52];
			partial_clause[448] 	= partial_clause_prev[448] & 1'b1;
			partial_clause[449] 	= partial_clause_prev[449] & 1'b1;
			partial_clause[450] 	= partial_clause_prev[450] & ~x[22] & ~x[23] & ~x[24] & ~x[26] & ~x[49];
			partial_clause[451] 	= partial_clause_prev[451] & 1'b1;
			partial_clause[452] 	= partial_clause_prev[452] & ~x[16] & ~x[21] & ~x[26];
			partial_clause[453] 	= partial_clause_prev[453] & ~x[20] & ~x[48];
			partial_clause[454] 	= partial_clause_prev[454] & ~x[2];
			partial_clause[455] 	= partial_clause_prev[455] & ~x[0] & ~x[1] & ~x[23] & ~x[51] & ~x[55];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[3] & ~x[23] & ~x[27] & ~x[28] & ~x[30] & ~x[52] & ~x[53] & ~x[56];
			partial_clause[457] 	= partial_clause_prev[457] & ~x[13] & ~x[14] & ~x[16] & ~x[37] & ~x[39] & ~x[47] & ~x[49];
			partial_clause[458] 	= partial_clause_prev[458] & ~x[17] & ~x[26] & ~x[45] & ~x[52] & ~x[53] & ~x[54] & ~x[58] & ~x[59];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[4] & ~x[6] & ~x[21] & ~x[32] & ~x[34] & ~x[48] & ~x[51] & ~x[53] & ~x[58] & ~x[59];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[2] & ~x[24] & ~x[30];
			partial_clause[461] 	= partial_clause_prev[461] & ~x[17] & ~x[25] & ~x[45];
			partial_clause[462] 	= partial_clause_prev[462] & ~x[32] & ~x[48];
			partial_clause[463] 	= partial_clause_prev[463] & ~x[51];
			partial_clause[464] 	= partial_clause_prev[464] & ~x[26] & ~x[53];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[22] & ~x[23] & ~x[24] & ~x[27] & ~x[28] & ~x[30] & ~x[52] & ~x[53] & ~x[57];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[0] & ~x[23] & ~x[24] & ~x[51] & ~x[55];
			partial_clause[467] 	= partial_clause_prev[467] & 1'b1;
			partial_clause[468] 	= partial_clause_prev[468] & ~x[0] & ~x[2] & ~x[21] & ~x[51];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[27];
			partial_clause[470] 	= partial_clause_prev[470] & 1'b1;
			partial_clause[471] 	= partial_clause_prev[471] & ~x[0] & ~x[4] & ~x[23] & ~x[28] & ~x[55] & ~x[59] & ~x[60];
			partial_clause[472] 	= partial_clause_prev[472] & x[42];
			partial_clause[473] 	= partial_clause_prev[473] & ~x[19] & ~x[23] & ~x[48];
			partial_clause[474] 	= partial_clause_prev[474] & ~x[2] & ~x[32] & ~x[48];
			partial_clause[475] 	= partial_clause_prev[475] & 1'b1;
			partial_clause[476] 	= partial_clause_prev[476] & 1'b1;
			partial_clause[477] 	= partial_clause_prev[477] & ~x[0] & ~x[21] & ~x[28] & ~x[50] & ~x[52] & ~x[53];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[16] & ~x[51] & ~x[53];
			partial_clause[479] 	= partial_clause_prev[479] & ~x[15] & ~x[16];
			partial_clause[480] 	= partial_clause_prev[480] & ~x[0] & ~x[20] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & ~x[46] & ~x[47] & ~x[49] & ~x[51] & ~x[52] & ~x[53] & ~x[55] & ~x[56];
			partial_clause[481] 	= partial_clause_prev[481] & ~x[27] & ~x[58];
			partial_clause[482] 	= partial_clause_prev[482] & ~x[24];
			partial_clause[483] 	= partial_clause_prev[483] & 1'b1;
			partial_clause[484] 	= partial_clause_prev[484] & ~x[35] & ~x[58] & ~x[63];
			partial_clause[485] 	= partial_clause_prev[485] & 1'b1;
			partial_clause[486] 	= partial_clause_prev[486] & ~x[1] & ~x[23];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[10] & ~x[27] & x[33] & ~x[55];
			partial_clause[488] 	= partial_clause_prev[488] & ~x[9] & ~x[37];
			partial_clause[489] 	= partial_clause_prev[489] & 1'b1;
			partial_clause[490] 	= partial_clause_prev[490] & ~x[7] & x[39];
			partial_clause[491] 	= partial_clause_prev[491] & ~x[51];
			partial_clause[492] 	= partial_clause_prev[492] & ~x[17] & ~x[18] & ~x[20] & ~x[53];
			partial_clause[493] 	= partial_clause_prev[493] & ~x[23];
			partial_clause[494] 	= partial_clause_prev[494] & ~x[22] & ~x[48] & ~x[53];
			partial_clause[495] 	= partial_clause_prev[495] & ~x[22] & ~x[50] & ~x[54];
			partial_clause[496] 	= partial_clause_prev[496] & 1'b1;
			partial_clause[497] 	= partial_clause_prev[497] & 1'b1;
			partial_clause[498] 	= partial_clause_prev[498] & 1'b1;
			partial_clause[499] 	= partial_clause_prev[499] & ~x[1] & ~x[12] & ~x[24] & ~x[40] & ~x[56];
		end
	end
endmodule


module HCB_5 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[13] & ~x[15] & ~x[17] & ~x[41] & ~x[44] & ~x[45] & ~x[49] & x[61];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[17] & ~x[21] & ~x[22] & ~x[37] & ~x[38] & ~x[49] & x[60];
			partial_clause[2] 	= partial_clause_prev[2] & ~x[11] & ~x[20];
			partial_clause[3] 	= partial_clause_prev[3] & 1'b1;
			partial_clause[4] 	= partial_clause_prev[4] & ~x[13] & ~x[20] & ~x[41] & ~x[58];
			partial_clause[5] 	= partial_clause_prev[5] & ~x[15] & ~x[18] & x[26] & ~x[42] & ~x[44] & ~x[47] & ~x[48] & ~x[50] & x[54];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[16] & ~x[18] & ~x[20] & ~x[40];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[16] & ~x[18] & ~x[21] & ~x[43] & ~x[44] & ~x[48];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[15] & ~x[20] & ~x[42] & ~x[45];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[16] & ~x[17] & ~x[43] & ~x[44] & ~x[47];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[14] & ~x[18] & ~x[43] & ~x[47] & x[63];
			partial_clause[11] 	= partial_clause_prev[11] & ~x[21] & ~x[40] & ~x[45] & ~x[50];
			partial_clause[12] 	= partial_clause_prev[12] & ~x[15] & ~x[18] & ~x[44] & ~x[46] & x[61];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[20] & ~x[21] & ~x[25] & ~x[46] & ~x[47] & ~x[50];
			partial_clause[14] 	= partial_clause_prev[14] & x[2] & ~x[22] & ~x[35];
			partial_clause[15] 	= partial_clause_prev[15] & 1'b1;
			partial_clause[16] 	= partial_clause_prev[16] & ~x[12] & ~x[38] & ~x[47];
			partial_clause[17] 	= partial_clause_prev[17] & x[57];
			partial_clause[18] 	= partial_clause_prev[18] & ~x[63];
			partial_clause[19] 	= partial_clause_prev[19] & ~x[10] & ~x[12] & ~x[37] & ~x[40];
			partial_clause[20] 	= partial_clause_prev[20] & ~x[57];
			partial_clause[21] 	= partial_clause_prev[21] & 1'b1;
			partial_clause[22] 	= partial_clause_prev[22] & ~x[3] & ~x[17] & ~x[58];
			partial_clause[23] 	= partial_clause_prev[23] & ~x[10] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[42] & ~x[43] & ~x[44] & ~x[45] & ~x[46] & ~x[47] & ~x[48] & ~x[49];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[15] & ~x[16] & ~x[17] & ~x[19] & ~x[20] & ~x[43] & ~x[44] & ~x[46] & ~x[49];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[14] & ~x[17] & ~x[22] & ~x[23] & ~x[38] & ~x[43] & ~x[44] & ~x[47] & ~x[49] & ~x[51];
			partial_clause[26] 	= partial_clause_prev[26] & x[56];
			partial_clause[27] 	= partial_clause_prev[27] & ~x[15] & ~x[21] & ~x[46] & ~x[48];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[46] & ~x[52];
			partial_clause[29] 	= partial_clause_prev[29] & x[6] & ~x[45] & x[60];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[22] & x[30] & ~x[38] & x[59];
			partial_clause[31] 	= partial_clause_prev[31] & 1'b1;
			partial_clause[32] 	= partial_clause_prev[32] & ~x[17] & ~x[53];
			partial_clause[33] 	= partial_clause_prev[33] & ~x[22];
			partial_clause[34] 	= partial_clause_prev[34] & ~x[45] & ~x[46] & ~x[47];
			partial_clause[35] 	= partial_clause_prev[35] & ~x[43] & ~x[44] & ~x[46];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[13] & ~x[51];
			partial_clause[37] 	= partial_clause_prev[37] & ~x[24];
			partial_clause[38] 	= partial_clause_prev[38] & ~x[9] & ~x[10] & ~x[15] & ~x[19] & ~x[41];
			partial_clause[39] 	= partial_clause_prev[39] & ~x[39] & ~x[52];
			partial_clause[40] 	= partial_clause_prev[40] & ~x[15] & ~x[19] & x[32] & ~x[39] & ~x[46] & x[58];
			partial_clause[41] 	= partial_clause_prev[41] & 1'b1;
			partial_clause[42] 	= partial_clause_prev[42] & ~x[1] & ~x[3] & ~x[26] & ~x[28] & ~x[52];
			partial_clause[43] 	= partial_clause_prev[43] & ~x[13] & ~x[18] & ~x[44] & ~x[46];
			partial_clause[44] 	= partial_clause_prev[44] & 1'b1;
			partial_clause[45] 	= partial_clause_prev[45] & x[32];
			partial_clause[46] 	= partial_clause_prev[46] & ~x[12] & ~x[16] & ~x[41] & ~x[47] & ~x[49];
			partial_clause[47] 	= partial_clause_prev[47] & ~x[18] & x[33] & ~x[38] & ~x[43];
			partial_clause[48] 	= partial_clause_prev[48] & 1'b1;
			partial_clause[49] 	= partial_clause_prev[49] & 1'b1;
			partial_clause[50] 	= partial_clause_prev[50] & ~x[3] & ~x[12] & ~x[40] & ~x[48];
			partial_clause[51] 	= partial_clause_prev[51] & 1'b1;
			partial_clause[52] 	= partial_clause_prev[52] & ~x[30];
			partial_clause[53] 	= partial_clause_prev[53] & ~x[4] & ~x[5] & ~x[6] & ~x[34] & ~x[35];
			partial_clause[54] 	= partial_clause_prev[54] & 1'b1;
			partial_clause[55] 	= partial_clause_prev[55] & ~x[4];
			partial_clause[56] 	= partial_clause_prev[56] & ~x[2];
			partial_clause[57] 	= partial_clause_prev[57] & ~x[11] & ~x[13] & ~x[19] & ~x[48];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[28];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[39] & ~x[40] & ~x[41] & ~x[44] & ~x[46];
			partial_clause[60] 	= partial_clause_prev[60] & 1'b1;
			partial_clause[61] 	= partial_clause_prev[61] & ~x[60];
			partial_clause[62] 	= partial_clause_prev[62] & ~x[12];
			partial_clause[63] 	= partial_clause_prev[63] & ~x[7] & ~x[32] & ~x[33];
			partial_clause[64] 	= partial_clause_prev[64] & ~x[1] & ~x[28] & ~x[43];
			partial_clause[65] 	= partial_clause_prev[65] & ~x[12] & ~x[26] & ~x[52];
			partial_clause[66] 	= partial_clause_prev[66] & x[10] & x[38];
			partial_clause[67] 	= partial_clause_prev[67] & x[31] & ~x[52];
			partial_clause[68] 	= partial_clause_prev[68] & 1'b1;
			partial_clause[69] 	= partial_clause_prev[69] & ~x[10] & ~x[13] & ~x[39] & ~x[40] & ~x[47];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[53] & ~x[54];
			partial_clause[71] 	= partial_clause_prev[71] & 1'b1;
			partial_clause[72] 	= partial_clause_prev[72] & x[7] & x[34];
			partial_clause[73] 	= partial_clause_prev[73] & ~x[28];
			partial_clause[74] 	= partial_clause_prev[74] & ~x[10] & ~x[18] & ~x[47];
			partial_clause[75] 	= partial_clause_prev[75] & 1'b1;
			partial_clause[76] 	= partial_clause_prev[76] & ~x[12] & ~x[19] & ~x[20] & ~x[41] & ~x[42] & ~x[47] & x[60];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[4];
			partial_clause[78] 	= partial_clause_prev[78] & ~x[9] & ~x[34] & ~x[46];
			partial_clause[79] 	= partial_clause_prev[79] & x[59];
			partial_clause[80] 	= partial_clause_prev[80] & ~x[2];
			partial_clause[81] 	= partial_clause_prev[81] & 1'b1;
			partial_clause[82] 	= partial_clause_prev[82] & ~x[42] & x[53];
			partial_clause[83] 	= partial_clause_prev[83] & ~x[0] & ~x[21];
			partial_clause[84] 	= partial_clause_prev[84] & 1'b1;
			partial_clause[85] 	= partial_clause_prev[85] & ~x[15] & ~x[21] & ~x[41] & ~x[43] & ~x[46] & ~x[50];
			partial_clause[86] 	= partial_clause_prev[86] & ~x[20] & ~x[39] & ~x[44];
			partial_clause[87] 	= partial_clause_prev[87] & ~x[15] & ~x[19] & ~x[36];
			partial_clause[88] 	= partial_clause_prev[88] & ~x[46] & ~x[47];
			partial_clause[89] 	= partial_clause_prev[89] & 1'b1;
			partial_clause[90] 	= partial_clause_prev[90] & 1'b1;
			partial_clause[91] 	= partial_clause_prev[91] & ~x[38] & x[60];
			partial_clause[92] 	= partial_clause_prev[92] & ~x[21] & ~x[43];
			partial_clause[93] 	= partial_clause_prev[93] & ~x[10] & ~x[11] & ~x[15] & ~x[17] & ~x[18] & ~x[38] & ~x[39] & ~x[44] & ~x[47] & ~x[48] & ~x[49];
			partial_clause[94] 	= partial_clause_prev[94] & 1'b1;
			partial_clause[95] 	= partial_clause_prev[95] & ~x[14] & ~x[35] & ~x[36] & ~x[63];
			partial_clause[96] 	= partial_clause_prev[96] & 1'b1;
			partial_clause[97] 	= partial_clause_prev[97] & ~x[19] & ~x[21] & ~x[38] & ~x[43] & x[55];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[15] & ~x[18] & ~x[20] & ~x[43] & ~x[45] & ~x[47] & ~x[48];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[12] & ~x[14] & ~x[15] & ~x[17] & ~x[28] & ~x[40] & ~x[41] & ~x[44] & ~x[45] & ~x[46] & ~x[47] & ~x[48];
			partial_clause[100] 	= partial_clause_prev[100] & ~x[11] & ~x[14] & ~x[41];
			partial_clause[101] 	= partial_clause_prev[101] & 1'b1;
			partial_clause[102] 	= partial_clause_prev[102] & ~x[17] & x[31] & ~x[39] & x[58];
			partial_clause[103] 	= partial_clause_prev[103] & ~x[10] & ~x[12] & ~x[13] & ~x[14] & ~x[16] & ~x[18] & ~x[21] & ~x[40] & ~x[49];
			partial_clause[104] 	= partial_clause_prev[104] & ~x[44];
			partial_clause[105] 	= partial_clause_prev[105] & ~x[13] & ~x[15] & ~x[17] & ~x[39];
			partial_clause[106] 	= partial_clause_prev[106] & ~x[44];
			partial_clause[107] 	= partial_clause_prev[107] & ~x[13] & ~x[20] & ~x[21] & ~x[39] & ~x[41] & ~x[47];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[11] & ~x[13] & ~x[15] & ~x[16] & ~x[20] & ~x[42] & ~x[45] & ~x[47];
			partial_clause[109] 	= partial_clause_prev[109] & 1'b1;
			partial_clause[110] 	= partial_clause_prev[110] & 1'b1;
			partial_clause[111] 	= partial_clause_prev[111] & x[23] & ~x[29];
			partial_clause[112] 	= partial_clause_prev[112] & ~x[43];
			partial_clause[113] 	= partial_clause_prev[113] & ~x[8] & ~x[19] & ~x[20];
			partial_clause[114] 	= partial_clause_prev[114] & 1'b1;
			partial_clause[115] 	= partial_clause_prev[115] & ~x[16] & ~x[22] & ~x[35] & ~x[36] & ~x[38] & ~x[43] & ~x[50];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[14] & ~x[15] & ~x[17] & ~x[18];
			partial_clause[117] 	= partial_clause_prev[117] & x[1] & ~x[7];
			partial_clause[118] 	= partial_clause_prev[118] & ~x[15] & ~x[18] & ~x[30] & ~x[41] & ~x[42] & ~x[45];
			partial_clause[119] 	= partial_clause_prev[119] & ~x[12] & ~x[15] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[47];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[14] & ~x[17] & ~x[43] & ~x[44] & ~x[46] & ~x[48];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[21] & ~x[23] & ~x[45];
			partial_clause[122] 	= partial_clause_prev[122] & ~x[43];
			partial_clause[123] 	= partial_clause_prev[123] & ~x[8] & ~x[9] & ~x[11] & ~x[17] & ~x[19] & ~x[39] & ~x[41] & ~x[42] & ~x[44] & ~x[45] & ~x[48] & ~x[50];
			partial_clause[124] 	= partial_clause_prev[124] & 1'b1;
			partial_clause[125] 	= partial_clause_prev[125] & ~x[15] & ~x[16] & ~x[47] & ~x[63];
			partial_clause[126] 	= partial_clause_prev[126] & 1'b1;
			partial_clause[127] 	= partial_clause_prev[127] & ~x[12] & ~x[19] & ~x[40] & ~x[42] & ~x[44] & ~x[46] & ~x[47] & ~x[48];
			partial_clause[128] 	= partial_clause_prev[128] & ~x[12] & ~x[13];
			partial_clause[129] 	= partial_clause_prev[129] & ~x[13] & ~x[16] & ~x[17] & ~x[40];
			partial_clause[130] 	= partial_clause_prev[130] & ~x[9] & ~x[16] & ~x[30] & ~x[49] & ~x[50];
			partial_clause[131] 	= partial_clause_prev[131] & 1'b1;
			partial_clause[132] 	= partial_clause_prev[132] & ~x[12] & ~x[46];
			partial_clause[133] 	= partial_clause_prev[133] & 1'b1;
			partial_clause[134] 	= partial_clause_prev[134] & ~x[15] & ~x[16] & ~x[37] & ~x[41] & ~x[43] & ~x[46] & ~x[47];
			partial_clause[135] 	= partial_clause_prev[135] & 1'b1;
			partial_clause[136] 	= partial_clause_prev[136] & ~x[12] & ~x[13] & ~x[40] & ~x[46];
			partial_clause[137] 	= partial_clause_prev[137] & x[63];
			partial_clause[138] 	= partial_clause_prev[138] & 1'b1;
			partial_clause[139] 	= partial_clause_prev[139] & ~x[10] & ~x[12] & ~x[13] & ~x[21] & ~x[36] & ~x[37] & ~x[38] & ~x[39] & ~x[40] & ~x[42] & ~x[45] & ~x[47];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[11] & ~x[15] & ~x[17] & ~x[41] & ~x[42] & ~x[45] & ~x[47] & ~x[51];
			partial_clause[141] 	= partial_clause_prev[141] & 1'b1;
			partial_clause[142] 	= partial_clause_prev[142] & ~x[47];
			partial_clause[143] 	= partial_clause_prev[143] & ~x[5] & x[8] & ~x[49];
			partial_clause[144] 	= partial_clause_prev[144] & ~x[36] & ~x[37] & ~x[38] & ~x[40] & x[54];
			partial_clause[145] 	= partial_clause_prev[145] & x[26] & x[55] & x[56];
			partial_clause[146] 	= partial_clause_prev[146] & 1'b1;
			partial_clause[147] 	= partial_clause_prev[147] & ~x[8] & ~x[13] & ~x[20] & ~x[39] & ~x[48] & ~x[49];
			partial_clause[148] 	= partial_clause_prev[148] & ~x[40] & ~x[42];
			partial_clause[149] 	= partial_clause_prev[149] & ~x[18] & ~x[47] & ~x[63];
			partial_clause[150] 	= partial_clause_prev[150] & ~x[11] & ~x[13] & ~x[26] & ~x[37] & ~x[38] & ~x[49] & ~x[53] & ~x[54];
			partial_clause[151] 	= partial_clause_prev[151] & ~x[54] & ~x[55];
			partial_clause[152] 	= partial_clause_prev[152] & 1'b1;
			partial_clause[153] 	= partial_clause_prev[153] & ~x[16] & ~x[17] & ~x[19] & ~x[41] & ~x[42] & ~x[43];
			partial_clause[154] 	= partial_clause_prev[154] & ~x[20];
			partial_clause[155] 	= partial_clause_prev[155] & 1'b1;
			partial_clause[156] 	= partial_clause_prev[156] & ~x[1] & ~x[19] & ~x[25] & ~x[26] & ~x[44];
			partial_clause[157] 	= partial_clause_prev[157] & 1'b1;
			partial_clause[158] 	= partial_clause_prev[158] & ~x[11] & ~x[15] & ~x[20] & ~x[41] & ~x[45] & ~x[46] & ~x[47] & x[61];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[11] & ~x[17] & ~x[19] & ~x[21] & ~x[22] & ~x[37] & ~x[39] & ~x[42] & ~x[49];
			partial_clause[160] 	= partial_clause_prev[160] & ~x[23];
			partial_clause[161] 	= partial_clause_prev[161] & ~x[12] & ~x[14] & ~x[16] & ~x[17] & ~x[38];
			partial_clause[162] 	= partial_clause_prev[162] & x[37];
			partial_clause[163] 	= partial_clause_prev[163] & ~x[60];
			partial_clause[164] 	= partial_clause_prev[164] & ~x[42] & ~x[47];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[11] & ~x[14] & ~x[16] & ~x[48];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[16] & ~x[42] & ~x[43] & ~x[45];
			partial_clause[167] 	= partial_clause_prev[167] & ~x[3];
			partial_clause[168] 	= partial_clause_prev[168] & ~x[11];
			partial_clause[169] 	= partial_clause_prev[169] & ~x[2] & ~x[18] & ~x[22] & ~x[29] & ~x[54] & ~x[55];
			partial_clause[170] 	= partial_clause_prev[170] & ~x[0];
			partial_clause[171] 	= partial_clause_prev[171] & ~x[12] & ~x[44] & x[52];
			partial_clause[172] 	= partial_clause_prev[172] & x[4];
			partial_clause[173] 	= partial_clause_prev[173] & ~x[11] & ~x[19] & ~x[41] & ~x[47];
			partial_clause[174] 	= partial_clause_prev[174] & ~x[13];
			partial_clause[175] 	= partial_clause_prev[175] & 1'b1;
			partial_clause[176] 	= partial_clause_prev[176] & ~x[18] & ~x[19] & ~x[21] & ~x[25] & ~x[28];
			partial_clause[177] 	= partial_clause_prev[177] & ~x[14] & ~x[40] & ~x[43];
			partial_clause[178] 	= partial_clause_prev[178] & 1'b1;
			partial_clause[179] 	= partial_clause_prev[179] & 1'b1;
			partial_clause[180] 	= partial_clause_prev[180] & ~x[45];
			partial_clause[181] 	= partial_clause_prev[181] & 1'b1;
			partial_clause[182] 	= partial_clause_prev[182] & 1'b1;
			partial_clause[183] 	= partial_clause_prev[183] & ~x[14] & ~x[17] & ~x[22] & ~x[37] & ~x[44] & ~x[50];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[47] & ~x[49];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[22];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[9] & ~x[16] & ~x[18] & ~x[20] & ~x[40] & ~x[46];
			partial_clause[187] 	= partial_clause_prev[187] & ~x[10] & ~x[11] & ~x[14] & ~x[15] & ~x[16] & ~x[41];
			partial_clause[188] 	= partial_clause_prev[188] & ~x[44];
			partial_clause[189] 	= partial_clause_prev[189] & 1'b1;
			partial_clause[190] 	= partial_clause_prev[190] & ~x[16] & x[61];
			partial_clause[191] 	= partial_clause_prev[191] & ~x[46];
			partial_clause[192] 	= partial_clause_prev[192] & ~x[8] & ~x[18] & ~x[20];
			partial_clause[193] 	= partial_clause_prev[193] & ~x[37] & ~x[47];
			partial_clause[194] 	= partial_clause_prev[194] & 1'b1;
			partial_clause[195] 	= partial_clause_prev[195] & ~x[13] & ~x[15] & ~x[43] & ~x[44];
			partial_clause[196] 	= partial_clause_prev[196] & 1'b1;
			partial_clause[197] 	= partial_clause_prev[197] & ~x[12] & ~x[19] & ~x[20] & ~x[24] & ~x[36] & ~x[43] & ~x[49];
			partial_clause[198] 	= partial_clause_prev[198] & 1'b1;
			partial_clause[199] 	= partial_clause_prev[199] & ~x[61];
			partial_clause[200] 	= partial_clause_prev[200] & ~x[11] & ~x[40];
			partial_clause[201] 	= partial_clause_prev[201] & ~x[14] & ~x[15] & ~x[41] & ~x[47] & ~x[50];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[10] & ~x[13] & ~x[16] & ~x[17] & ~x[19] & ~x[21] & ~x[40] & ~x[41] & ~x[43] & ~x[44] & ~x[46];
			partial_clause[203] 	= partial_clause_prev[203] & ~x[12] & ~x[27] & ~x[53];
			partial_clause[204] 	= partial_clause_prev[204] & ~x[42] & ~x[45] & ~x[47];
			partial_clause[205] 	= partial_clause_prev[205] & 1'b1;
			partial_clause[206] 	= partial_clause_prev[206] & ~x[13] & ~x[14] & ~x[16] & ~x[44] & ~x[47];
			partial_clause[207] 	= partial_clause_prev[207] & ~x[16] & ~x[21] & ~x[39] & ~x[46];
			partial_clause[208] 	= partial_clause_prev[208] & x[33] & ~x[43] & x[61];
			partial_clause[209] 	= partial_clause_prev[209] & ~x[9];
			partial_clause[210] 	= partial_clause_prev[210] & ~x[10] & ~x[12] & ~x[22] & ~x[41] & ~x[43] & ~x[50];
			partial_clause[211] 	= partial_clause_prev[211] & 1'b1;
			partial_clause[212] 	= partial_clause_prev[212] & ~x[11] & ~x[14] & ~x[21] & ~x[47];
			partial_clause[213] 	= partial_clause_prev[213] & 1'b1;
			partial_clause[214] 	= partial_clause_prev[214] & ~x[50];
			partial_clause[215] 	= partial_clause_prev[215] & ~x[20];
			partial_clause[216] 	= partial_clause_prev[216] & 1'b1;
			partial_clause[217] 	= partial_clause_prev[217] & ~x[13] & ~x[44];
			partial_clause[218] 	= partial_clause_prev[218] & ~x[33] & ~x[34] & ~x[61];
			partial_clause[219] 	= partial_clause_prev[219] & 1'b1;
			partial_clause[220] 	= partial_clause_prev[220] & 1'b1;
			partial_clause[221] 	= partial_clause_prev[221] & ~x[16] & ~x[39] & ~x[57];
			partial_clause[222] 	= partial_clause_prev[222] & x[54];
			partial_clause[223] 	= partial_clause_prev[223] & ~x[14];
			partial_clause[224] 	= partial_clause_prev[224] & ~x[12] & ~x[16] & ~x[37] & ~x[41] & ~x[42] & ~x[49];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[16] & x[31] & ~x[38];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[16] & ~x[18] & ~x[44] & ~x[45] & ~x[46];
			partial_clause[227] 	= partial_clause_prev[227] & ~x[18];
			partial_clause[228] 	= partial_clause_prev[228] & ~x[23] & ~x[44] & ~x[50];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[16] & ~x[40] & ~x[41] & ~x[46] & ~x[48];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[15] & ~x[19] & ~x[21] & ~x[38] & ~x[39] & ~x[42] & ~x[49] & ~x[50] & x[55];
			partial_clause[231] 	= partial_clause_prev[231] & ~x[13] & ~x[20] & ~x[32] & ~x[44] & ~x[48];
			partial_clause[232] 	= partial_clause_prev[232] & ~x[32] & ~x[60];
			partial_clause[233] 	= partial_clause_prev[233] & 1'b1;
			partial_clause[234] 	= partial_clause_prev[234] & ~x[13] & ~x[25] & ~x[29] & ~x[44];
			partial_clause[235] 	= partial_clause_prev[235] & ~x[2] & ~x[30];
			partial_clause[236] 	= partial_clause_prev[236] & ~x[53];
			partial_clause[237] 	= partial_clause_prev[237] & 1'b1;
			partial_clause[238] 	= partial_clause_prev[238] & 1'b1;
			partial_clause[239] 	= partial_clause_prev[239] & 1'b1;
			partial_clause[240] 	= partial_clause_prev[240] & ~x[38] & ~x[41] & ~x[44];
			partial_clause[241] 	= partial_clause_prev[241] & x[62];
			partial_clause[242] 	= partial_clause_prev[242] & ~x[13] & ~x[14] & ~x[17] & ~x[21] & ~x[42] & ~x[45] & ~x[46] & ~x[47] & ~x[48];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[1] & ~x[47] & ~x[48] & ~x[54] & ~x[55];
			partial_clause[244] 	= partial_clause_prev[244] & ~x[1] & ~x[13] & ~x[43];
			partial_clause[245] 	= partial_clause_prev[245] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[11] & ~x[34] & ~x[35] & ~x[37];
			partial_clause[246] 	= partial_clause_prev[246] & ~x[53] & x[57];
			partial_clause[247] 	= partial_clause_prev[247] & ~x[12] & ~x[21] & ~x[41] & ~x[45] & ~x[47];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[11] & ~x[15] & ~x[19] & ~x[20] & ~x[42] & ~x[44] & ~x[47] & ~x[48];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[6] & ~x[10] & ~x[14] & ~x[16] & ~x[36] & ~x[38] & ~x[39];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[15] & ~x[20] & ~x[40] & ~x[43] & ~x[46] & ~x[49] & ~x[50];
			partial_clause[251] 	= partial_clause_prev[251] & ~x[12];
			partial_clause[252] 	= partial_clause_prev[252] & ~x[15] & ~x[19] & ~x[20] & ~x[22] & ~x[37] & ~x[41] & ~x[44] & ~x[50];
			partial_clause[253] 	= partial_clause_prev[253] & ~x[9] & ~x[21] & ~x[23] & ~x[41];
			partial_clause[254] 	= partial_clause_prev[254] & ~x[2] & ~x[19];
			partial_clause[255] 	= partial_clause_prev[255] & ~x[13] & ~x[17] & ~x[19] & ~x[20];
			partial_clause[256] 	= partial_clause_prev[256] & x[26];
			partial_clause[257] 	= partial_clause_prev[257] & ~x[2];
			partial_clause[258] 	= partial_clause_prev[258] & ~x[2] & ~x[40] & ~x[43] & ~x[46];
			partial_clause[259] 	= partial_clause_prev[259] & 1'b1;
			partial_clause[260] 	= partial_clause_prev[260] & ~x[12] & ~x[39];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[23] & ~x[48];
			partial_clause[262] 	= partial_clause_prev[262] & ~x[19] & ~x[48];
			partial_clause[263] 	= partial_clause_prev[263] & 1'b1;
			partial_clause[264] 	= partial_clause_prev[264] & ~x[39] & ~x[46];
			partial_clause[265] 	= partial_clause_prev[265] & 1'b1;
			partial_clause[266] 	= partial_clause_prev[266] & ~x[11] & ~x[13] & ~x[20] & ~x[22] & ~x[39] & ~x[40] & ~x[41] & ~x[43];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[19] & ~x[20] & ~x[40] & ~x[41] & ~x[42] & ~x[44] & ~x[48];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[14] & ~x[21] & x[27];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[14] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[42] & ~x[45] & ~x[46];
			partial_clause[270] 	= partial_clause_prev[270] & x[30];
			partial_clause[271] 	= partial_clause_prev[271] & 1'b1;
			partial_clause[272] 	= partial_clause_prev[272] & ~x[18] & ~x[20] & x[33] & ~x[44] & ~x[45];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[11] & ~x[12] & ~x[14] & ~x[15] & ~x[17] & ~x[18] & ~x[19] & ~x[41];
			partial_clause[274] 	= partial_clause_prev[274] & ~x[16] & ~x[19] & ~x[21];
			partial_clause[275] 	= partial_clause_prev[275] & 1'b1;
			partial_clause[276] 	= partial_clause_prev[276] & ~x[10] & x[59];
			partial_clause[277] 	= partial_clause_prev[277] & ~x[4] & ~x[40];
			partial_clause[278] 	= partial_clause_prev[278] & 1'b1;
			partial_clause[279] 	= partial_clause_prev[279] & ~x[9] & ~x[12] & ~x[17] & ~x[20] & ~x[22] & ~x[37] & ~x[39] & ~x[40] & ~x[45] & ~x[48] & ~x[49];
			partial_clause[280] 	= partial_clause_prev[280] & x[25];
			partial_clause[281] 	= partial_clause_prev[281] & ~x[18] & ~x[19] & ~x[41] & ~x[47];
			partial_clause[282] 	= partial_clause_prev[282] & ~x[13] & ~x[14] & ~x[45];
			partial_clause[283] 	= partial_clause_prev[283] & 1'b1;
			partial_clause[284] 	= partial_clause_prev[284] & x[31] & ~x[36] & ~x[48];
			partial_clause[285] 	= partial_clause_prev[285] & ~x[51];
			partial_clause[286] 	= partial_clause_prev[286] & ~x[40] & ~x[45];
			partial_clause[287] 	= partial_clause_prev[287] & ~x[11] & ~x[18] & ~x[20] & ~x[22] & ~x[38] & ~x[39] & ~x[51];
			partial_clause[288] 	= partial_clause_prev[288] & 1'b1;
			partial_clause[289] 	= partial_clause_prev[289] & ~x[39] & ~x[44];
			partial_clause[290] 	= partial_clause_prev[290] & ~x[18] & ~x[41];
			partial_clause[291] 	= partial_clause_prev[291] & 1'b1;
			partial_clause[292] 	= partial_clause_prev[292] & ~x[18] & ~x[46];
			partial_clause[293] 	= partial_clause_prev[293] & x[6] & ~x[13] & ~x[14] & ~x[29];
			partial_clause[294] 	= partial_clause_prev[294] & ~x[12] & ~x[46];
			partial_clause[295] 	= partial_clause_prev[295] & ~x[1] & ~x[28] & ~x[29] & ~x[44] & ~x[55];
			partial_clause[296] 	= partial_clause_prev[296] & x[5] & ~x[16] & ~x[22] & ~x[57] & ~x[58];
			partial_clause[297] 	= partial_clause_prev[297] & ~x[13];
			partial_clause[298] 	= partial_clause_prev[298] & 1'b1;
			partial_clause[299] 	= partial_clause_prev[299] & ~x[17] & ~x[39];
			partial_clause[300] 	= partial_clause_prev[300] & ~x[24] & ~x[41] & ~x[43];
			partial_clause[301] 	= partial_clause_prev[301] & ~x[49];
			partial_clause[302] 	= partial_clause_prev[302] & ~x[10] & ~x[17] & ~x[44];
			partial_clause[303] 	= partial_clause_prev[303] & ~x[30];
			partial_clause[304] 	= partial_clause_prev[304] & ~x[12] & ~x[15] & ~x[17] & ~x[47];
			partial_clause[305] 	= partial_clause_prev[305] & 1'b1;
			partial_clause[306] 	= partial_clause_prev[306] & ~x[15] & ~x[19] & ~x[48];
			partial_clause[307] 	= partial_clause_prev[307] & ~x[10] & ~x[22] & ~x[38] & ~x[47] & ~x[50];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[47] & ~x[54];
			partial_clause[309] 	= partial_clause_prev[309] & ~x[16] & ~x[31] & ~x[41] & ~x[44] & ~x[58];
			partial_clause[310] 	= partial_clause_prev[310] & ~x[3] & ~x[5] & ~x[7] & ~x[8] & ~x[36];
			partial_clause[311] 	= partial_clause_prev[311] & 1'b1;
			partial_clause[312] 	= partial_clause_prev[312] & x[54];
			partial_clause[313] 	= partial_clause_prev[313] & ~x[12] & ~x[17] & ~x[40];
			partial_clause[314] 	= partial_clause_prev[314] & ~x[43];
			partial_clause[315] 	= partial_clause_prev[315] & ~x[12];
			partial_clause[316] 	= partial_clause_prev[316] & ~x[14] & ~x[22] & ~x[37] & ~x[41] & ~x[44] & ~x[45] & ~x[46];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[11] & ~x[16] & ~x[43];
			partial_clause[318] 	= partial_clause_prev[318] & ~x[6] & ~x[10] & ~x[35] & ~x[40] & ~x[42] & ~x[48];
			partial_clause[319] 	= partial_clause_prev[319] & ~x[17] & ~x[35] & ~x[44] & ~x[62] & ~x[63];
			partial_clause[320] 	= partial_clause_prev[320] & ~x[15] & ~x[18] & ~x[20] & ~x[43] & ~x[48] & ~x[50] & ~x[52] & ~x[53] & ~x[54];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[12] & ~x[18] & ~x[19] & ~x[20] & ~x[22] & ~x[41] & ~x[42] & ~x[45];
			partial_clause[322] 	= partial_clause_prev[322] & ~x[19] & ~x[21] & ~x[45];
			partial_clause[323] 	= partial_clause_prev[323] & 1'b1;
			partial_clause[324] 	= partial_clause_prev[324] & ~x[34] & ~x[48];
			partial_clause[325] 	= partial_clause_prev[325] & ~x[13] & ~x[14] & ~x[16] & ~x[19] & ~x[21] & ~x[22] & ~x[23] & ~x[40] & ~x[43] & ~x[48];
			partial_clause[326] 	= partial_clause_prev[326] & x[23] & ~x[43] & ~x[44] & ~x[45] & ~x[46];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[11] & ~x[15] & ~x[50];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[19] & ~x[24] & ~x[28] & ~x[48] & ~x[52] & ~x[55];
			partial_clause[329] 	= partial_clause_prev[329] & x[34];
			partial_clause[330] 	= partial_clause_prev[330] & ~x[13] & ~x[46];
			partial_clause[331] 	= partial_clause_prev[331] & ~x[14] & x[33] & x[34] & ~x[48] & x[59];
			partial_clause[332] 	= partial_clause_prev[332] & ~x[1] & ~x[2] & ~x[18] & ~x[19];
			partial_clause[333] 	= partial_clause_prev[333] & ~x[0] & ~x[22] & ~x[23];
			partial_clause[334] 	= partial_clause_prev[334] & x[0] & ~x[9] & ~x[14] & ~x[20] & ~x[38] & ~x[41];
			partial_clause[335] 	= partial_clause_prev[335] & 1'b1;
			partial_clause[336] 	= partial_clause_prev[336] & x[3];
			partial_clause[337] 	= partial_clause_prev[337] & ~x[13] & ~x[25] & ~x[41] & ~x[46] & ~x[48];
			partial_clause[338] 	= partial_clause_prev[338] & 1'b1;
			partial_clause[339] 	= partial_clause_prev[339] & ~x[10] & ~x[20] & ~x[40] & ~x[47] & ~x[50];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[14] & ~x[16] & ~x[17] & ~x[40] & ~x[43] & ~x[45] & ~x[46];
			partial_clause[341] 	= partial_clause_prev[341] & x[57];
			partial_clause[342] 	= partial_clause_prev[342] & ~x[11] & ~x[12] & ~x[13] & ~x[16] & ~x[37] & ~x[47] & ~x[48];
			partial_clause[343] 	= partial_clause_prev[343] & ~x[11] & ~x[12] & ~x[14] & ~x[18] & ~x[19];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[6] & ~x[12] & ~x[15] & ~x[18] & ~x[23] & ~x[47];
			partial_clause[345] 	= partial_clause_prev[345] & x[28] & ~x[37];
			partial_clause[346] 	= partial_clause_prev[346] & ~x[17] & ~x[29] & ~x[57];
			partial_clause[347] 	= partial_clause_prev[347] & 1'b1;
			partial_clause[348] 	= partial_clause_prev[348] & 1'b1;
			partial_clause[349] 	= partial_clause_prev[349] & ~x[16] & ~x[31] & ~x[45];
			partial_clause[350] 	= partial_clause_prev[350] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[42] & ~x[44] & x[60];
			partial_clause[351] 	= partial_clause_prev[351] & ~x[4];
			partial_clause[352] 	= partial_clause_prev[352] & x[10];
			partial_clause[353] 	= partial_clause_prev[353] & ~x[57];
			partial_clause[354] 	= partial_clause_prev[354] & ~x[13] & ~x[17] & ~x[44];
			partial_clause[355] 	= partial_clause_prev[355] & ~x[17] & ~x[41];
			partial_clause[356] 	= partial_clause_prev[356] & 1'b1;
			partial_clause[357] 	= partial_clause_prev[357] & 1'b1;
			partial_clause[358] 	= partial_clause_prev[358] & ~x[15] & ~x[46];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[17] & ~x[40];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[13] & ~x[16] & ~x[17];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[14] & ~x[44];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[45];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[10] & ~x[11] & ~x[12] & ~x[22] & ~x[37] & ~x[39] & ~x[43] & ~x[47];
			partial_clause[364] 	= partial_clause_prev[364] & ~x[12] & ~x[21];
			partial_clause[365] 	= partial_clause_prev[365] & 1'b1;
			partial_clause[366] 	= partial_clause_prev[366] & ~x[42] & ~x[45] & ~x[47] & x[61];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[21] & ~x[40] & ~x[47];
			partial_clause[368] 	= partial_clause_prev[368] & 1'b1;
			partial_clause[369] 	= partial_clause_prev[369] & ~x[14] & ~x[40];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[10] & ~x[37] & ~x[39] & ~x[49];
			partial_clause[371] 	= partial_clause_prev[371] & 1'b1;
			partial_clause[372] 	= partial_clause_prev[372] & x[5];
			partial_clause[373] 	= partial_clause_prev[373] & 1'b1;
			partial_clause[374] 	= partial_clause_prev[374] & ~x[19] & ~x[20];
			partial_clause[375] 	= partial_clause_prev[375] & ~x[27] & ~x[50] & ~x[52];
			partial_clause[376] 	= partial_clause_prev[376] & ~x[9] & ~x[15] & ~x[17] & ~x[22];
			partial_clause[377] 	= partial_clause_prev[377] & ~x[46];
			partial_clause[378] 	= partial_clause_prev[378] & ~x[37] & ~x[40] & ~x[50];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[0] & ~x[1] & ~x[25] & ~x[52];
			partial_clause[380] 	= partial_clause_prev[380] & ~x[39];
			partial_clause[381] 	= partial_clause_prev[381] & ~x[13] & ~x[14] & ~x[41] & ~x[43] & ~x[49];
			partial_clause[382] 	= partial_clause_prev[382] & ~x[5] & ~x[32];
			partial_clause[383] 	= partial_clause_prev[383] & ~x[41] & x[58];
			partial_clause[384] 	= partial_clause_prev[384] & 1'b1;
			partial_clause[385] 	= partial_clause_prev[385] & 1'b1;
			partial_clause[386] 	= partial_clause_prev[386] & ~x[17] & ~x[59];
			partial_clause[387] 	= partial_clause_prev[387] & ~x[10] & ~x[12] & ~x[14] & ~x[16] & ~x[18] & ~x[19] & ~x[21] & ~x[22] & ~x[39] & ~x[44] & ~x[50] & ~x[63];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[3] & ~x[16] & ~x[17] & ~x[18] & ~x[44] & ~x[45];
			partial_clause[389] 	= partial_clause_prev[389] & 1'b1;
			partial_clause[390] 	= partial_clause_prev[390] & ~x[11] & ~x[48];
			partial_clause[391] 	= partial_clause_prev[391] & 1'b1;
			partial_clause[392] 	= partial_clause_prev[392] & 1'b1;
			partial_clause[393] 	= partial_clause_prev[393] & x[3];
			partial_clause[394] 	= partial_clause_prev[394] & ~x[18] & ~x[22] & ~x[38];
			partial_clause[395] 	= partial_clause_prev[395] & ~x[20];
			partial_clause[396] 	= partial_clause_prev[396] & ~x[49];
			partial_clause[397] 	= partial_clause_prev[397] & ~x[27] & ~x[45];
			partial_clause[398] 	= partial_clause_prev[398] & ~x[7] & ~x[37];
			partial_clause[399] 	= partial_clause_prev[399] & 1'b1;
			partial_clause[400] 	= partial_clause_prev[400] & ~x[17] & ~x[39] & ~x[45];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[11] & ~x[15] & ~x[21] & ~x[38] & ~x[39] & ~x[44] & ~x[47] & ~x[48] & ~x[50];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[38] & ~x[44] & ~x[45] & x[59];
			partial_clause[403] 	= partial_clause_prev[403] & 1'b1;
			partial_clause[404] 	= partial_clause_prev[404] & 1'b1;
			partial_clause[405] 	= partial_clause_prev[405] & ~x[18] & ~x[42] & ~x[46];
			partial_clause[406] 	= partial_clause_prev[406] & ~x[7] & ~x[12] & ~x[24] & ~x[49];
			partial_clause[407] 	= partial_clause_prev[407] & ~x[8] & x[27] & ~x[39] & ~x[46];
			partial_clause[408] 	= partial_clause_prev[408] & ~x[40] & ~x[44] & ~x[47];
			partial_clause[409] 	= partial_clause_prev[409] & ~x[9] & ~x[16] & ~x[17] & ~x[18] & ~x[20] & ~x[21] & ~x[22] & ~x[43] & ~x[45] & ~x[49] & ~x[50];
			partial_clause[410] 	= partial_clause_prev[410] & ~x[8] & ~x[46];
			partial_clause[411] 	= partial_clause_prev[411] & ~x[10] & ~x[15] & ~x[16];
			partial_clause[412] 	= partial_clause_prev[412] & ~x[10] & ~x[13] & ~x[16] & ~x[21] & ~x[35] & ~x[36] & ~x[44] & ~x[46] & ~x[49] & ~x[62];
			partial_clause[413] 	= partial_clause_prev[413] & ~x[13];
			partial_clause[414] 	= partial_clause_prev[414] & ~x[16] & ~x[18] & ~x[21] & ~x[22] & ~x[44] & ~x[46] & ~x[48];
			partial_clause[415] 	= partial_clause_prev[415] & ~x[6] & ~x[21] & ~x[23] & ~x[40] & ~x[45] & ~x[46] & ~x[47] & ~x[50];
			partial_clause[416] 	= partial_clause_prev[416] & ~x[16] & ~x[19] & ~x[24] & ~x[44] & ~x[49];
			partial_clause[417] 	= partial_clause_prev[417] & ~x[15];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[10] & ~x[11] & ~x[14] & ~x[16] & ~x[20] & ~x[22] & ~x[38] & ~x[40] & ~x[42] & ~x[43] & ~x[44] & ~x[45] & ~x[47];
			partial_clause[419] 	= partial_clause_prev[419] & ~x[22];
			partial_clause[420] 	= partial_clause_prev[420] & ~x[26];
			partial_clause[421] 	= partial_clause_prev[421] & ~x[30] & ~x[42];
			partial_clause[422] 	= partial_clause_prev[422] & ~x[14] & ~x[27] & ~x[46];
			partial_clause[423] 	= partial_clause_prev[423] & ~x[11] & ~x[20] & ~x[45] & ~x[47] & ~x[50];
			partial_clause[424] 	= partial_clause_prev[424] & ~x[41] & x[59];
			partial_clause[425] 	= partial_clause_prev[425] & 1'b1;
			partial_clause[426] 	= partial_clause_prev[426] & ~x[20] & ~x[44] & ~x[46] & ~x[47];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[17] & ~x[36] & ~x[40] & ~x[42] & ~x[43] & ~x[44];
			partial_clause[428] 	= partial_clause_prev[428] & 1'b1;
			partial_clause[429] 	= partial_clause_prev[429] & ~x[24];
			partial_clause[430] 	= partial_clause_prev[430] & ~x[13] & ~x[18] & ~x[19] & ~x[45] & ~x[51];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[15] & ~x[20] & ~x[38] & x[58] & x[59];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[11] & ~x[15] & ~x[17] & ~x[19] & ~x[22] & ~x[40] & ~x[46] & ~x[48] & ~x[49] & ~x[50];
			partial_clause[433] 	= partial_clause_prev[433] & ~x[13] & ~x[17] & ~x[19] & ~x[45];
			partial_clause[434] 	= partial_clause_prev[434] & 1'b1;
			partial_clause[435] 	= partial_clause_prev[435] & ~x[12] & ~x[14] & ~x[16] & ~x[17] & ~x[18] & x[33] & ~x[50] & ~x[52];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[12] & ~x[15] & ~x[17] & ~x[18] & ~x[21] & ~x[23] & ~x[41] & ~x[47];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[14] & ~x[19] & ~x[20] & ~x[22] & ~x[45] & ~x[49];
			partial_clause[438] 	= partial_clause_prev[438] & 1'b1;
			partial_clause[439] 	= partial_clause_prev[439] & ~x[10] & ~x[16] & ~x[22] & ~x[37] & ~x[39] & ~x[42] & ~x[47] & ~x[48] & ~x[50];
			partial_clause[440] 	= partial_clause_prev[440] & ~x[21];
			partial_clause[441] 	= partial_clause_prev[441] & x[28];
			partial_clause[442] 	= partial_clause_prev[442] & ~x[57];
			partial_clause[443] 	= partial_clause_prev[443] & ~x[11] & ~x[14] & ~x[18] & ~x[19] & ~x[44] & x[59] & x[60];
			partial_clause[444] 	= partial_clause_prev[444] & ~x[59];
			partial_clause[445] 	= partial_clause_prev[445] & ~x[43] & ~x[57];
			partial_clause[446] 	= partial_clause_prev[446] & ~x[41] & ~x[45] & ~x[47];
			partial_clause[447] 	= partial_clause_prev[447] & ~x[13] & ~x[44];
			partial_clause[448] 	= partial_clause_prev[448] & 1'b1;
			partial_clause[449] 	= partial_clause_prev[449] & ~x[15] & ~x[18] & x[28] & ~x[36] & ~x[45] & ~x[49];
			partial_clause[450] 	= partial_clause_prev[450] & 1'b1;
			partial_clause[451] 	= partial_clause_prev[451] & ~x[25];
			partial_clause[452] 	= partial_clause_prev[452] & ~x[8] & ~x[37];
			partial_clause[453] 	= partial_clause_prev[453] & ~x[42];
			partial_clause[454] 	= partial_clause_prev[454] & ~x[16];
			partial_clause[455] 	= partial_clause_prev[455] & ~x[44] & x[59];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[47] & ~x[48];
			partial_clause[457] 	= partial_clause_prev[457] & 1'b1;
			partial_clause[458] 	= partial_clause_prev[458] & ~x[9] & ~x[17] & ~x[19] & ~x[20] & x[30] & ~x[40] & ~x[41] & ~x[50];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[21] & ~x[40] & ~x[43] & ~x[44] & ~x[45];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[6] & ~x[11] & ~x[12] & ~x[35];
			partial_clause[461] 	= partial_clause_prev[461] & ~x[18];
			partial_clause[462] 	= partial_clause_prev[462] & ~x[36] & ~x[40];
			partial_clause[463] 	= partial_clause_prev[463] & ~x[28] & ~x[54];
			partial_clause[464] 	= partial_clause_prev[464] & ~x[12];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[16] & ~x[48] & ~x[50];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[13] & ~x[14] & ~x[15] & ~x[43] & ~x[46];
			partial_clause[467] 	= partial_clause_prev[467] & ~x[10];
			partial_clause[468] 	= partial_clause_prev[468] & ~x[22] & ~x[42];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[55];
			partial_clause[470] 	= partial_clause_prev[470] & ~x[0] & ~x[38] & ~x[53] & ~x[54];
			partial_clause[471] 	= partial_clause_prev[471] & ~x[11] & ~x[40] & ~x[41] & ~x[45] & ~x[46];
			partial_clause[472] 	= partial_clause_prev[472] & ~x[23];
			partial_clause[473] 	= partial_clause_prev[473] & ~x[11] & ~x[13] & ~x[15] & ~x[20] & ~x[22] & ~x[41] & ~x[45];
			partial_clause[474] 	= partial_clause_prev[474] & 1'b1;
			partial_clause[475] 	= partial_clause_prev[475] & ~x[14];
			partial_clause[476] 	= partial_clause_prev[476] & 1'b1;
			partial_clause[477] 	= partial_clause_prev[477] & ~x[2] & ~x[12] & ~x[18] & ~x[22] & ~x[24] & ~x[25] & ~x[28] & ~x[29] & ~x[45];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[13] & ~x[39];
			partial_clause[479] 	= partial_clause_prev[479] & 1'b1;
			partial_clause[480] 	= partial_clause_prev[480] & ~x[12] & ~x[13] & ~x[16] & ~x[18] & ~x[19] & ~x[21] & ~x[22] & ~x[38] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[47] & ~x[48] & ~x[49] & ~x[50];
			partial_clause[481] 	= partial_clause_prev[481] & ~x[28] & ~x[51];
			partial_clause[482] 	= partial_clause_prev[482] & ~x[2] & ~x[41] & ~x[43] & ~x[55];
			partial_clause[483] 	= partial_clause_prev[483] & ~x[35] & x[57];
			partial_clause[484] 	= partial_clause_prev[484] & ~x[20] & ~x[22];
			partial_clause[485] 	= partial_clause_prev[485] & 1'b1;
			partial_clause[486] 	= partial_clause_prev[486] & ~x[3] & ~x[13] & ~x[16] & ~x[30] & ~x[45];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[15] & ~x[20] & ~x[42];
			partial_clause[488] 	= partial_clause_prev[488] & 1'b1;
			partial_clause[489] 	= partial_clause_prev[489] & 1'b1;
			partial_clause[490] 	= partial_clause_prev[490] & 1'b1;
			partial_clause[491] 	= partial_clause_prev[491] & ~x[2] & x[60];
			partial_clause[492] 	= partial_clause_prev[492] & ~x[13] & ~x[14] & ~x[16] & ~x[43];
			partial_clause[493] 	= partial_clause_prev[493] & ~x[18] & ~x[28] & ~x[38] & ~x[52] & ~x[54];
			partial_clause[494] 	= partial_clause_prev[494] & ~x[40];
			partial_clause[495] 	= partial_clause_prev[495] & ~x[11] & ~x[19] & ~x[20] & ~x[42] & ~x[45];
			partial_clause[496] 	= partial_clause_prev[496] & 1'b1;
			partial_clause[497] 	= partial_clause_prev[497] & ~x[56];
			partial_clause[498] 	= partial_clause_prev[498] & ~x[19] & ~x[59];
			partial_clause[499] 	= partial_clause_prev[499] & ~x[2] & ~x[13];
		end
	end
endmodule


module HCB_6 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[6] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & x[22] & x[23] & ~x[32] & ~x[34] & ~x[36] & ~x[38] & x[50] & ~x[61] & ~x[62];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[13] & ~x[34] & ~x[38] & ~x[43] & ~x[56];
			partial_clause[2] 	= partial_clause_prev[2] & ~x[37];
			partial_clause[3] 	= partial_clause_prev[3] & ~x[2] & ~x[29];
			partial_clause[4] 	= partial_clause_prev[4] & x[44];
			partial_clause[5] 	= partial_clause_prev[5] & ~x[8] & ~x[9] & ~x[12] & ~x[14] & x[18] & ~x[35] & ~x[40] & ~x[41] & ~x[61];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[10] & ~x[36] & ~x[38] & ~x[40];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[0] & ~x[10] & ~x[25] & ~x[26] & ~x[30] & ~x[40] & ~x[55];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[2] & ~x[4] & ~x[6] & ~x[9] & ~x[11] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[37];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[8] & ~x[10] & ~x[30] & ~x[33] & ~x[34];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[4] & ~x[8] & ~x[33] & ~x[39] & ~x[42];
			partial_clause[11] 	= partial_clause_prev[11] & ~x[12] & ~x[13] & ~x[33] & ~x[36] & ~x[38] & ~x[40];
			partial_clause[12] 	= partial_clause_prev[12] & ~x[7] & ~x[9] & ~x[33] & ~x[35] & ~x[37];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[6] & ~x[7] & ~x[11] & ~x[14] & ~x[15] & ~x[30] & ~x[38] & ~x[41] & ~x[55] & ~x[56] & ~x[59];
			partial_clause[14] 	= partial_clause_prev[14] & ~x[2] & ~x[3] & ~x[43];
			partial_clause[15] 	= partial_clause_prev[15] & ~x[20] & ~x[40];
			partial_clause[16] 	= partial_clause_prev[16] & ~x[10] & x[26] & ~x[31] & x[53] & ~x[57] & ~x[58] & ~x[60] & ~x[62];
			partial_clause[17] 	= partial_clause_prev[17] & ~x[41];
			partial_clause[18] 	= partial_clause_prev[18] & ~x[0] & ~x[61];
			partial_clause[19] 	= partial_clause_prev[19] & ~x[2] & ~x[34] & ~x[35] & ~x[39] & ~x[61];
			partial_clause[20] 	= partial_clause_prev[20] & 1'b1;
			partial_clause[21] 	= partial_clause_prev[21] & 1'b1;
			partial_clause[22] 	= partial_clause_prev[22] & ~x[31] & ~x[34];
			partial_clause[23] 	= partial_clause_prev[23] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[12] & ~x[13] & ~x[33] & ~x[34] & ~x[36] & ~x[37] & ~x[38] & ~x[39] & ~x[40] & ~x[62] & ~x[63];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[6] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[33] & ~x[34] & ~x[36] & ~x[37] & ~x[38] & ~x[39] & ~x[40] & ~x[62];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[1] & ~x[2] & ~x[6] & ~x[8] & ~x[10] & ~x[12] & ~x[37] & ~x[39] & ~x[40] & ~x[41] & ~x[57] & ~x[62];
			partial_clause[26] 	= partial_clause_prev[26] & 1'b1;
			partial_clause[27] 	= partial_clause_prev[27] & ~x[5];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[7] & ~x[14] & ~x[27] & ~x[28] & ~x[36] & ~x[43];
			partial_clause[29] 	= partial_clause_prev[29] & ~x[30] & x[49] & x[50] & ~x[57];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[15] & ~x[33] & ~x[35] & ~x[41] & ~x[60] & ~x[61];
			partial_clause[31] 	= partial_clause_prev[31] & ~x[42] & ~x[63];
			partial_clause[32] 	= partial_clause_prev[32] & ~x[15] & ~x[17] & ~x[32] & ~x[43] & ~x[59];
			partial_clause[33] 	= partial_clause_prev[33] & ~x[31];
			partial_clause[34] 	= partial_clause_prev[34] & ~x[8] & ~x[11] & ~x[34] & ~x[39];
			partial_clause[35] 	= partial_clause_prev[35] & ~x[6] & ~x[7] & ~x[32] & ~x[35] & ~x[38];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[8] & ~x[9] & ~x[13] & ~x[20] & ~x[31] & ~x[43] & ~x[45];
			partial_clause[37] 	= partial_clause_prev[37] & x[20] & ~x[40];
			partial_clause[38] 	= partial_clause_prev[38] & ~x[9] & ~x[31] & ~x[34];
			partial_clause[39] 	= partial_clause_prev[39] & ~x[13] & ~x[16];
			partial_clause[40] 	= partial_clause_prev[40] & ~x[10] & ~x[36] & ~x[61];
			partial_clause[41] 	= partial_clause_prev[41] & x[46];
			partial_clause[42] 	= partial_clause_prev[42] & ~x[3] & ~x[42];
			partial_clause[43] 	= partial_clause_prev[43] & ~x[34] & ~x[38] & x[50] & ~x[63];
			partial_clause[44] 	= partial_clause_prev[44] & ~x[48];
			partial_clause[45] 	= partial_clause_prev[45] & ~x[7] & x[23];
			partial_clause[46] 	= partial_clause_prev[46] & ~x[2] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[29] & ~x[32] & ~x[34] & ~x[35] & ~x[38] & ~x[39] & ~x[42] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[47] 	= partial_clause_prev[47] & ~x[4] & ~x[12] & x[53] & ~x[61];
			partial_clause[48] 	= partial_clause_prev[48] & 1'b1;
			partial_clause[49] 	= partial_clause_prev[49] & ~x[31] & ~x[38];
			partial_clause[50] 	= partial_clause_prev[50] & ~x[37] & ~x[41];
			partial_clause[51] 	= partial_clause_prev[51] & x[15] & ~x[20];
			partial_clause[52] 	= partial_clause_prev[52] & x[1];
			partial_clause[53] 	= partial_clause_prev[53] & ~x[2] & ~x[59];
			partial_clause[54] 	= partial_clause_prev[54] & x[27] & x[55];
			partial_clause[55] 	= partial_clause_prev[55] & 1'b1;
			partial_clause[56] 	= partial_clause_prev[56] & 1'b1;
			partial_clause[57] 	= partial_clause_prev[57] & ~x[36];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[11] & ~x[16] & ~x[17] & ~x[31] & ~x[33] & ~x[40] & ~x[60];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[3] & ~x[4] & ~x[32] & ~x[35] & ~x[38] & ~x[62];
			partial_clause[60] 	= partial_clause_prev[60] & 1'b1;
			partial_clause[61] 	= partial_clause_prev[61] & ~x[42] & ~x[52];
			partial_clause[62] 	= partial_clause_prev[62] & ~x[11] & ~x[60] & ~x[62];
			partial_clause[63] 	= partial_clause_prev[63] & ~x[10] & ~x[38];
			partial_clause[64] 	= partial_clause_prev[64] & ~x[3];
			partial_clause[65] 	= partial_clause_prev[65] & ~x[14] & x[49] & x[50];
			partial_clause[66] 	= partial_clause_prev[66] & 1'b1;
			partial_clause[67] 	= partial_clause_prev[67] & 1'b1;
			partial_clause[68] 	= partial_clause_prev[68] & ~x[37] & ~x[46] & ~x[49];
			partial_clause[69] 	= partial_clause_prev[69] & ~x[12] & ~x[29] & ~x[35] & ~x[40] & x[51];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[33] & ~x[36] & ~x[59] & ~x[60];
			partial_clause[71] 	= partial_clause_prev[71] & ~x[9] & ~x[13] & x[23] & ~x[43] & ~x[61] & ~x[63];
			partial_clause[72] 	= partial_clause_prev[72] & 1'b1;
			partial_clause[73] 	= partial_clause_prev[73] & 1'b1;
			partial_clause[74] 	= partial_clause_prev[74] & ~x[7] & ~x[11] & ~x[39] & ~x[42] & ~x[43];
			partial_clause[75] 	= partial_clause_prev[75] & ~x[19] & ~x[47];
			partial_clause[76] 	= partial_clause_prev[76] & ~x[1] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[10] & ~x[12] & ~x[14] & ~x[32] & ~x[34] & ~x[40] & ~x[60] & ~x[62];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[5] & ~x[60];
			partial_clause[78] 	= partial_clause_prev[78] & ~x[24];
			partial_clause[79] 	= partial_clause_prev[79] & ~x[5];
			partial_clause[80] 	= partial_clause_prev[80] & 1'b1;
			partial_clause[81] 	= partial_clause_prev[81] & ~x[13] & ~x[34];
			partial_clause[82] 	= partial_clause_prev[82] & x[44];
			partial_clause[83] 	= partial_clause_prev[83] & ~x[56];
			partial_clause[84] 	= partial_clause_prev[84] & 1'b1;
			partial_clause[85] 	= partial_clause_prev[85] & ~x[5] & ~x[32] & ~x[34] & ~x[42] & ~x[62] & ~x[63];
			partial_clause[86] 	= partial_clause_prev[86] & ~x[39];
			partial_clause[87] 	= partial_clause_prev[87] & ~x[2] & ~x[39];
			partial_clause[88] 	= partial_clause_prev[88] & ~x[50];
			partial_clause[89] 	= partial_clause_prev[89] & ~x[46] & ~x[47];
			partial_clause[90] 	= partial_clause_prev[90] & ~x[3];
			partial_clause[91] 	= partial_clause_prev[91] & ~x[8] & ~x[32] & ~x[58];
			partial_clause[92] 	= partial_clause_prev[92] & ~x[3] & ~x[36] & ~x[37] & ~x[41] & ~x[59];
			partial_clause[93] 	= partial_clause_prev[93] & ~x[1] & ~x[4] & ~x[5] & ~x[10] & ~x[11] & ~x[15] & ~x[31] & ~x[33] & ~x[34] & ~x[35] & ~x[37] & ~x[38] & ~x[58];
			partial_clause[94] 	= partial_clause_prev[94] & ~x[22];
			partial_clause[95] 	= partial_clause_prev[95] & ~x[7] & ~x[9] & ~x[11] & ~x[36] & ~x[57] & ~x[63];
			partial_clause[96] 	= partial_clause_prev[96] & ~x[48] & ~x[49] & ~x[50];
			partial_clause[97] 	= partial_clause_prev[97] & ~x[4] & ~x[6] & ~x[8] & ~x[9] & ~x[13] & ~x[14] & ~x[39] & ~x[42] & ~x[43] & ~x[44] & ~x[58] & ~x[60];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[7] & ~x[9] & ~x[12] & ~x[40] & ~x[61];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[2] & ~x[3] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[31] & ~x[32] & ~x[33] & ~x[35] & ~x[38] & ~x[57] & ~x[58] & ~x[59] & ~x[60] & ~x[63];
			partial_clause[100] 	= partial_clause_prev[100] & 1'b1;
			partial_clause[101] 	= partial_clause_prev[101] & x[19] & x[21];
			partial_clause[102] 	= partial_clause_prev[102] & ~x[0];
			partial_clause[103] 	= partial_clause_prev[103] & ~x[1] & ~x[4] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[12] & ~x[20] & ~x[36] & ~x[38] & ~x[39] & ~x[40] & ~x[41] & ~x[43] & ~x[59] & ~x[63];
			partial_clause[104] 	= partial_clause_prev[104] & ~x[33];
			partial_clause[105] 	= partial_clause_prev[105] & ~x[6] & ~x[9] & ~x[34] & ~x[38] & ~x[41];
			partial_clause[106] 	= partial_clause_prev[106] & ~x[8] & ~x[12] & ~x[59] & ~x[60];
			partial_clause[107] 	= partial_clause_prev[107] & ~x[35] & ~x[39] & ~x[40] & x[52] & ~x[61] & ~x[62];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[8] & ~x[32] & ~x[33] & ~x[61] & ~x[63];
			partial_clause[109] 	= partial_clause_prev[109] & 1'b1;
			partial_clause[110] 	= partial_clause_prev[110] & 1'b1;
			partial_clause[111] 	= partial_clause_prev[111] & x[14];
			partial_clause[112] 	= partial_clause_prev[112] & ~x[9] & ~x[34];
			partial_clause[113] 	= partial_clause_prev[113] & ~x[10] & x[53];
			partial_clause[114] 	= partial_clause_prev[114] & 1'b1;
			partial_clause[115] 	= partial_clause_prev[115] & ~x[1] & ~x[4] & ~x[7] & ~x[8] & ~x[12] & ~x[13] & ~x[32] & ~x[36] & ~x[41] & ~x[43] & ~x[62];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[3] & ~x[36] & ~x[39] & ~x[58] & ~x[61];
			partial_clause[117] 	= partial_clause_prev[117] & 1'b1;
			partial_clause[118] 	= partial_clause_prev[118] & ~x[13] & ~x[35];
			partial_clause[119] 	= partial_clause_prev[119] & ~x[5] & ~x[6] & ~x[7] & ~x[12] & ~x[36] & ~x[38] & ~x[40];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[3] & ~x[7] & ~x[9] & ~x[12] & ~x[33] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[39] & ~x[40] & ~x[60] & ~x[62];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[5] & ~x[32] & ~x[34] & ~x[39] & ~x[61];
			partial_clause[122] 	= partial_clause_prev[122] & ~x[7] & ~x[13] & ~x[14] & ~x[26] & ~x[34] & ~x[55] & ~x[61];
			partial_clause[123] 	= partial_clause_prev[123] & ~x[2] & ~x[8] & ~x[11] & ~x[12] & ~x[13] & ~x[32] & ~x[33] & ~x[36] & ~x[37] & ~x[39] & ~x[41] & ~x[59];
			partial_clause[124] 	= partial_clause_prev[124] & 1'b1;
			partial_clause[125] 	= partial_clause_prev[125] & ~x[5] & ~x[29] & ~x[54];
			partial_clause[126] 	= partial_clause_prev[126] & x[22] & x[23];
			partial_clause[127] 	= partial_clause_prev[127] & ~x[5] & ~x[7] & ~x[12] & ~x[33] & ~x[44] & ~x[62];
			partial_clause[128] 	= partial_clause_prev[128] & ~x[5] & ~x[9] & ~x[31] & ~x[32] & ~x[63];
			partial_clause[129] 	= partial_clause_prev[129] & ~x[9] & ~x[13] & ~x[36] & ~x[38] & ~x[58] & ~x[60] & ~x[61];
			partial_clause[130] 	= partial_clause_prev[130] & ~x[7] & ~x[21];
			partial_clause[131] 	= partial_clause_prev[131] & ~x[32] & ~x[33];
			partial_clause[132] 	= partial_clause_prev[132] & ~x[7] & ~x[35] & ~x[37];
			partial_clause[133] 	= partial_clause_prev[133] & ~x[7] & x[52];
			partial_clause[134] 	= partial_clause_prev[134] & ~x[0] & ~x[1] & ~x[2] & ~x[6] & ~x[10] & x[20] & ~x[31] & ~x[32] & ~x[34] & ~x[35] & ~x[37] & ~x[40] & ~x[57] & ~x[63];
			partial_clause[135] 	= partial_clause_prev[135] & 1'b1;
			partial_clause[136] 	= partial_clause_prev[136] & ~x[3] & ~x[5] & ~x[12] & ~x[37] & ~x[42] & ~x[63];
			partial_clause[137] 	= partial_clause_prev[137] & ~x[31] & x[53];
			partial_clause[138] 	= partial_clause_prev[138] & 1'b1;
			partial_clause[139] 	= partial_clause_prev[139] & ~x[0] & ~x[1] & ~x[6] & ~x[7] & ~x[9] & x[22] & ~x[28] & ~x[29] & ~x[30] & ~x[38] & ~x[41];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[0] & ~x[13] & ~x[15] & ~x[31] & ~x[32] & ~x[33] & ~x[34] & ~x[43] & ~x[58] & ~x[60];
			partial_clause[141] 	= partial_clause_prev[141] & ~x[34];
			partial_clause[142] 	= partial_clause_prev[142] & ~x[6] & ~x[33] & ~x[36];
			partial_clause[143] 	= partial_clause_prev[143] & ~x[31] & ~x[58] & ~x[60] & ~x[61];
			partial_clause[144] 	= partial_clause_prev[144] & ~x[11] & ~x[63];
			partial_clause[145] 	= partial_clause_prev[145] & 1'b1;
			partial_clause[146] 	= partial_clause_prev[146] & ~x[36] & x[49] & x[50];
			partial_clause[147] 	= partial_clause_prev[147] & ~x[9] & ~x[14] & ~x[34];
			partial_clause[148] 	= partial_clause_prev[148] & ~x[5] & ~x[7];
			partial_clause[149] 	= partial_clause_prev[149] & ~x[27] & ~x[30] & ~x[58];
			partial_clause[150] 	= partial_clause_prev[150] & ~x[2] & ~x[9] & ~x[18] & ~x[29] & ~x[35] & ~x[38] & ~x[40];
			partial_clause[151] 	= partial_clause_prev[151] & 1'b1;
			partial_clause[152] 	= partial_clause_prev[152] & 1'b1;
			partial_clause[153] 	= partial_clause_prev[153] & ~x[36] & ~x[37] & ~x[38] & ~x[63];
			partial_clause[154] 	= partial_clause_prev[154] & x[22] & x[49] & ~x[54];
			partial_clause[155] 	= partial_clause_prev[155] & 1'b1;
			partial_clause[156] 	= partial_clause_prev[156] & ~x[16];
			partial_clause[157] 	= partial_clause_prev[157] & x[3];
			partial_clause[158] 	= partial_clause_prev[158] & ~x[1] & ~x[6] & ~x[7] & ~x[11] & ~x[31] & ~x[37] & ~x[39] & ~x[41] & ~x[55] & ~x[57];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[2] & ~x[27] & ~x[35] & ~x[54] & ~x[58] & ~x[63];
			partial_clause[160] 	= partial_clause_prev[160] & ~x[8] & ~x[12] & ~x[16] & ~x[27] & ~x[55] & ~x[56];
			partial_clause[161] 	= partial_clause_prev[161] & ~x[6] & ~x[9] & ~x[10] & ~x[14] & ~x[42] & ~x[61];
			partial_clause[162] 	= partial_clause_prev[162] & ~x[6] & ~x[11] & ~x[37] & ~x[63];
			partial_clause[163] 	= partial_clause_prev[163] & 1'b1;
			partial_clause[164] 	= partial_clause_prev[164] & ~x[4] & ~x[6] & ~x[44];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[38];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[6] & ~x[37];
			partial_clause[167] 	= partial_clause_prev[167] & 1'b1;
			partial_clause[168] 	= partial_clause_prev[168] & ~x[1] & ~x[30] & ~x[32] & ~x[33] & ~x[63];
			partial_clause[169] 	= partial_clause_prev[169] & ~x[8] & ~x[16] & ~x[43];
			partial_clause[170] 	= partial_clause_prev[170] & 1'b1;
			partial_clause[171] 	= partial_clause_prev[171] & ~x[10] & ~x[12] & ~x[32] & ~x[38];
			partial_clause[172] 	= partial_clause_prev[172] & 1'b1;
			partial_clause[173] 	= partial_clause_prev[173] & ~x[3] & ~x[5] & ~x[9] & ~x[38] & ~x[60];
			partial_clause[174] 	= partial_clause_prev[174] & x[23] & x[24];
			partial_clause[175] 	= partial_clause_prev[175] & 1'b1;
			partial_clause[176] 	= partial_clause_prev[176] & ~x[6] & ~x[61];
			partial_clause[177] 	= partial_clause_prev[177] & ~x[37];
			partial_clause[178] 	= partial_clause_prev[178] & x[25] & ~x[40] & x[52] & ~x[57];
			partial_clause[179] 	= partial_clause_prev[179] & 1'b1;
			partial_clause[180] 	= partial_clause_prev[180] & 1'b1;
			partial_clause[181] 	= partial_clause_prev[181] & 1'b1;
			partial_clause[182] 	= partial_clause_prev[182] & x[54];
			partial_clause[183] 	= partial_clause_prev[183] & ~x[14] & ~x[33] & ~x[43] & ~x[61];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[4] & ~x[6] & ~x[12] & ~x[29] & ~x[34] & ~x[58];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[5];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[4] & ~x[9] & ~x[33] & ~x[37] & ~x[39] & ~x[55];
			partial_clause[187] 	= partial_clause_prev[187] & ~x[5] & ~x[8] & ~x[11] & ~x[34] & ~x[36] & ~x[38] & ~x[59];
			partial_clause[188] 	= partial_clause_prev[188] & ~x[38];
			partial_clause[189] 	= partial_clause_prev[189] & ~x[22];
			partial_clause[190] 	= partial_clause_prev[190] & ~x[35] & ~x[60] & ~x[63];
			partial_clause[191] 	= partial_clause_prev[191] & ~x[44];
			partial_clause[192] 	= partial_clause_prev[192] & ~x[10];
			partial_clause[193] 	= partial_clause_prev[193] & ~x[8] & ~x[29] & ~x[55] & ~x[57] & ~x[60] & ~x[62];
			partial_clause[194] 	= partial_clause_prev[194] & 1'b1;
			partial_clause[195] 	= partial_clause_prev[195] & ~x[2] & ~x[13] & ~x[29] & ~x[31] & ~x[33] & ~x[36] & ~x[56] & ~x[61];
			partial_clause[196] 	= partial_clause_prev[196] & 1'b1;
			partial_clause[197] 	= partial_clause_prev[197] & ~x[4] & ~x[14] & ~x[35] & ~x[36] & ~x[37] & ~x[40];
			partial_clause[198] 	= partial_clause_prev[198] & ~x[1];
			partial_clause[199] 	= partial_clause_prev[199] & 1'b1;
			partial_clause[200] 	= partial_clause_prev[200] & ~x[9] & ~x[34] & ~x[35];
			partial_clause[201] 	= partial_clause_prev[201] & ~x[4] & ~x[39] & ~x[41];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[4] & ~x[7] & ~x[9] & ~x[10] & ~x[12] & ~x[16] & ~x[33] & ~x[39] & ~x[41] & ~x[60] & ~x[63];
			partial_clause[203] 	= partial_clause_prev[203] & ~x[4] & ~x[16] & ~x[35] & ~x[41] & x[49];
			partial_clause[204] 	= partial_clause_prev[204] & ~x[10] & ~x[33] & ~x[36];
			partial_clause[205] 	= partial_clause_prev[205] & 1'b1;
			partial_clause[206] 	= partial_clause_prev[206] & ~x[4] & ~x[15] & x[21] & x[22] & ~x[36] & ~x[38] & ~x[59];
			partial_clause[207] 	= partial_clause_prev[207] & ~x[8] & ~x[11] & ~x[16] & ~x[30] & ~x[32] & ~x[59] & ~x[60];
			partial_clause[208] 	= partial_clause_prev[208] & ~x[37] & ~x[61];
			partial_clause[209] 	= partial_clause_prev[209] & 1'b1;
			partial_clause[210] 	= partial_clause_prev[210] & ~x[2] & ~x[4] & ~x[10] & ~x[11] & ~x[35] & ~x[36] & ~x[38] & ~x[40] & ~x[58] & ~x[59];
			partial_clause[211] 	= partial_clause_prev[211] & ~x[0] & ~x[26] & ~x[54];
			partial_clause[212] 	= partial_clause_prev[212] & ~x[42] & ~x[61];
			partial_clause[213] 	= partial_clause_prev[213] & 1'b1;
			partial_clause[214] 	= partial_clause_prev[214] & ~x[41];
			partial_clause[215] 	= partial_clause_prev[215] & 1'b1;
			partial_clause[216] 	= partial_clause_prev[216] & ~x[9] & ~x[44];
			partial_clause[217] 	= partial_clause_prev[217] & ~x[22] & ~x[37] & ~x[63];
			partial_clause[218] 	= partial_clause_prev[218] & ~x[36];
			partial_clause[219] 	= partial_clause_prev[219] & ~x[39];
			partial_clause[220] 	= partial_clause_prev[220] & ~x[33] & ~x[34] & ~x[58];
			partial_clause[221] 	= partial_clause_prev[221] & ~x[12];
			partial_clause[222] 	= partial_clause_prev[222] & x[17] & x[45] & x[46];
			partial_clause[223] 	= partial_clause_prev[223] & ~x[31] & ~x[41] & x[51];
			partial_clause[224] 	= partial_clause_prev[224] & ~x[2] & ~x[33] & ~x[39] & ~x[60];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[37] & ~x[40] & ~x[60];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[4] & ~x[5] & ~x[7] & ~x[9] & ~x[30] & ~x[33] & ~x[34] & ~x[36] & ~x[60] & ~x[63];
			partial_clause[227] 	= partial_clause_prev[227] & 1'b1;
			partial_clause[228] 	= partial_clause_prev[228] & ~x[5] & ~x[8] & ~x[12] & ~x[28] & ~x[29] & ~x[35] & ~x[40] & ~x[58] & ~x[62];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[10] & ~x[13] & ~x[31] & ~x[36] & ~x[37] & ~x[55] & ~x[58] & ~x[62] & ~x[63];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[1] & ~x[4] & ~x[6] & ~x[9] & ~x[11] & ~x[12] & ~x[13] & x[19] & ~x[28] & ~x[32] & ~x[35] & ~x[37] & ~x[40] & ~x[59] & ~x[60] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[231] 	= partial_clause_prev[231] & ~x[11];
			partial_clause[232] 	= partial_clause_prev[232] & ~x[24] & ~x[51];
			partial_clause[233] 	= partial_clause_prev[233] & ~x[59];
			partial_clause[234] 	= partial_clause_prev[234] & 1'b1;
			partial_clause[235] 	= partial_clause_prev[235] & ~x[21];
			partial_clause[236] 	= partial_clause_prev[236] & ~x[11] & ~x[15];
			partial_clause[237] 	= partial_clause_prev[237] & ~x[7] & ~x[31] & ~x[39];
			partial_clause[238] 	= partial_clause_prev[238] & ~x[56];
			partial_clause[239] 	= partial_clause_prev[239] & ~x[17] & x[51];
			partial_clause[240] 	= partial_clause_prev[240] & ~x[2] & ~x[11] & ~x[12] & ~x[29];
			partial_clause[241] 	= partial_clause_prev[241] & x[26] & ~x[30] & ~x[32] & ~x[59];
			partial_clause[242] 	= partial_clause_prev[242] & ~x[4] & ~x[9] & x[19] & ~x[39] & ~x[40] & ~x[61];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[12] & ~x[18];
			partial_clause[244] 	= partial_clause_prev[244] & 1'b1;
			partial_clause[245] 	= partial_clause_prev[245] & ~x[33];
			partial_clause[246] 	= partial_clause_prev[246] & ~x[5] & ~x[32] & ~x[43];
			partial_clause[247] 	= partial_clause_prev[247] & ~x[4] & ~x[6] & ~x[7] & ~x[12] & ~x[13] & ~x[32] & ~x[41] & ~x[42] & ~x[62] & ~x[63];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[3] & ~x[5] & ~x[8] & ~x[13] & ~x[31] & ~x[32] & ~x[40] & ~x[42] & ~x[61] & ~x[63];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[31] & ~x[34];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[3] & ~x[4] & ~x[6] & ~x[7] & ~x[8] & ~x[12] & ~x[13] & ~x[14] & ~x[29] & ~x[31] & ~x[32] & ~x[34] & ~x[37] & ~x[38] & ~x[40] & ~x[41] & ~x[42] & ~x[44] & ~x[56] & ~x[59] & ~x[61];
			partial_clause[251] 	= partial_clause_prev[251] & ~x[42];
			partial_clause[252] 	= partial_clause_prev[252] & ~x[15] & ~x[16] & ~x[33] & ~x[34] & ~x[36] & ~x[60];
			partial_clause[253] 	= partial_clause_prev[253] & ~x[5] & ~x[10];
			partial_clause[254] 	= partial_clause_prev[254] & ~x[8] & ~x[11] & ~x[31] & ~x[60];
			partial_clause[255] 	= partial_clause_prev[255] & ~x[9] & ~x[11];
			partial_clause[256] 	= partial_clause_prev[256] & 1'b1;
			partial_clause[257] 	= partial_clause_prev[257] & x[23] & x[24] & ~x[32] & x[49];
			partial_clause[258] 	= partial_clause_prev[258] & ~x[5] & x[45] & ~x[62];
			partial_clause[259] 	= partial_clause_prev[259] & x[15] & x[30] & x[43];
			partial_clause[260] 	= partial_clause_prev[260] & ~x[2] & ~x[19] & ~x[20] & ~x[47] & ~x[48] & ~x[63];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[7] & ~x[12] & ~x[32] & ~x[34] & ~x[44];
			partial_clause[262] 	= partial_clause_prev[262] & 1'b1;
			partial_clause[263] 	= partial_clause_prev[263] & 1'b1;
			partial_clause[264] 	= partial_clause_prev[264] & ~x[11] & x[23] & ~x[35] & ~x[57] & ~x[62];
			partial_clause[265] 	= partial_clause_prev[265] & ~x[45];
			partial_clause[266] 	= partial_clause_prev[266] & ~x[1] & ~x[4] & ~x[63];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[8] & ~x[10] & ~x[36] & ~x[37] & ~x[38] & ~x[61];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[6] & ~x[9] & ~x[29] & ~x[31] & ~x[36] & ~x[37] & ~x[40] & ~x[59] & ~x[62];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[6] & ~x[8] & ~x[9] & ~x[12] & ~x[33] & ~x[34] & ~x[35] & ~x[36] & ~x[38] & ~x[60] & ~x[61] & ~x[63];
			partial_clause[270] 	= partial_clause_prev[270] & x[22];
			partial_clause[271] 	= partial_clause_prev[271] & ~x[20];
			partial_clause[272] 	= partial_clause_prev[272] & ~x[8] & ~x[11] & ~x[36] & ~x[37] & x[48];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[5] & ~x[8] & ~x[10] & ~x[32] & ~x[33] & ~x[36] & ~x[38] & ~x[39] & ~x[40] & ~x[62];
			partial_clause[274] 	= partial_clause_prev[274] & ~x[37] & ~x[38] & ~x[62];
			partial_clause[275] 	= partial_clause_prev[275] & ~x[5];
			partial_clause[276] 	= partial_clause_prev[276] & ~x[2] & x[23] & ~x[33] & ~x[43];
			partial_clause[277] 	= partial_clause_prev[277] & ~x[4] & ~x[13];
			partial_clause[278] 	= partial_clause_prev[278] & ~x[24];
			partial_clause[279] 	= partial_clause_prev[279] & ~x[0] & ~x[28] & ~x[29] & ~x[36] & ~x[40] & ~x[58] & ~x[61];
			partial_clause[280] 	= partial_clause_prev[280] & x[16];
			partial_clause[281] 	= partial_clause_prev[281] & ~x[14] & ~x[33] & ~x[36];
			partial_clause[282] 	= partial_clause_prev[282] & ~x[6] & ~x[12] & ~x[39] & ~x[62];
			partial_clause[283] 	= partial_clause_prev[283] & x[51];
			partial_clause[284] 	= partial_clause_prev[284] & ~x[0] & ~x[8] & ~x[54];
			partial_clause[285] 	= partial_clause_prev[285] & ~x[9] & ~x[13];
			partial_clause[286] 	= partial_clause_prev[286] & ~x[35] & ~x[36];
			partial_clause[287] 	= partial_clause_prev[287] & ~x[0] & ~x[1] & ~x[2] & ~x[4] & ~x[5] & ~x[8] & ~x[9] & ~x[15] & ~x[28] & ~x[30] & ~x[31] & ~x[32] & ~x[38] & ~x[39] & ~x[40] & ~x[59] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[288] 	= partial_clause_prev[288] & ~x[21] & ~x[37];
			partial_clause[289] 	= partial_clause_prev[289] & ~x[41];
			partial_clause[290] 	= partial_clause_prev[290] & ~x[11] & ~x[14] & ~x[15] & ~x[58];
			partial_clause[291] 	= partial_clause_prev[291] & 1'b1;
			partial_clause[292] 	= partial_clause_prev[292] & ~x[13] & ~x[37] & ~x[40];
			partial_clause[293] 	= partial_clause_prev[293] & ~x[58];
			partial_clause[294] 	= partial_clause_prev[294] & ~x[6] & x[24] & ~x[31] & ~x[38] & ~x[39] & x[52];
			partial_clause[295] 	= partial_clause_prev[295] & ~x[8] & ~x[13] & ~x[15] & ~x[17];
			partial_clause[296] 	= partial_clause_prev[296] & 1'b1;
			partial_clause[297] 	= partial_clause_prev[297] & ~x[31] & ~x[58];
			partial_clause[298] 	= partial_clause_prev[298] & 1'b1;
			partial_clause[299] 	= partial_clause_prev[299] & ~x[3] & ~x[10] & ~x[59];
			partial_clause[300] 	= partial_clause_prev[300] & ~x[38] & ~x[41];
			partial_clause[301] 	= partial_clause_prev[301] & ~x[7] & ~x[35] & ~x[37] & ~x[39] & ~x[61];
			partial_clause[302] 	= partial_clause_prev[302] & ~x[5] & ~x[63];
			partial_clause[303] 	= partial_clause_prev[303] & ~x[14];
			partial_clause[304] 	= partial_clause_prev[304] & 1'b1;
			partial_clause[305] 	= partial_clause_prev[305] & ~x[11] & ~x[38] & ~x[41];
			partial_clause[306] 	= partial_clause_prev[306] & 1'b1;
			partial_clause[307] 	= partial_clause_prev[307] & ~x[2] & ~x[4] & ~x[42] & ~x[43] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[15] & ~x[29] & ~x[33] & ~x[39] & ~x[61] & ~x[62];
			partial_clause[309] 	= partial_clause_prev[309] & ~x[8] & ~x[22] & ~x[35] & ~x[49] & ~x[50] & ~x[61];
			partial_clause[310] 	= partial_clause_prev[310] & ~x[1] & ~x[2];
			partial_clause[311] 	= partial_clause_prev[311] & ~x[8];
			partial_clause[312] 	= partial_clause_prev[312] & ~x[23] & ~x[62];
			partial_clause[313] 	= partial_clause_prev[313] & 1'b1;
			partial_clause[314] 	= partial_clause_prev[314] & ~x[6] & ~x[36] & ~x[39];
			partial_clause[315] 	= partial_clause_prev[315] & ~x[33];
			partial_clause[316] 	= partial_clause_prev[316] & ~x[7] & ~x[8] & ~x[30] & ~x[31] & ~x[36] & ~x[38] & ~x[39] & ~x[41] & ~x[56] & ~x[59] & ~x[60] & ~x[61];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[3] & ~x[32];
			partial_clause[318] 	= partial_clause_prev[318] & ~x[1] & ~x[30] & ~x[38];
			partial_clause[319] 	= partial_clause_prev[319] & ~x[38] & ~x[63];
			partial_clause[320] 	= partial_clause_prev[320] & ~x[8] & ~x[9] & ~x[13] & ~x[14] & ~x[63];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[3] & ~x[5] & ~x[11] & ~x[12] & ~x[15] & ~x[16] & x[21] & ~x[34] & ~x[40] & x[50] & ~x[57] & ~x[60];
			partial_clause[322] 	= partial_clause_prev[322] & ~x[4] & ~x[7] & ~x[14] & ~x[43] & ~x[58];
			partial_clause[323] 	= partial_clause_prev[323] & ~x[4] & ~x[5] & ~x[11];
			partial_clause[324] 	= partial_clause_prev[324] & 1'b1;
			partial_clause[325] 	= partial_clause_prev[325] & ~x[3] & ~x[10] & ~x[13] & ~x[32] & ~x[35] & ~x[37] & ~x[38] & ~x[39] & ~x[40] & ~x[59] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[326] 	= partial_clause_prev[326] & ~x[6] & ~x[9];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[14] & ~x[31] & ~x[34] & ~x[61];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[34] & ~x[35] & ~x[40] & ~x[61];
			partial_clause[329] 	= partial_clause_prev[329] & ~x[35];
			partial_clause[330] 	= partial_clause_prev[330] & ~x[7] & ~x[31] & x[49];
			partial_clause[331] 	= partial_clause_prev[331] & ~x[4] & x[22] & ~x[29] & ~x[31] & ~x[57] & ~x[58] & ~x[62];
			partial_clause[332] 	= partial_clause_prev[332] & ~x[10] & ~x[11] & ~x[39] & ~x[58];
			partial_clause[333] 	= partial_clause_prev[333] & 1'b1;
			partial_clause[334] 	= partial_clause_prev[334] & ~x[4] & ~x[6] & ~x[38] & ~x[62];
			partial_clause[335] 	= partial_clause_prev[335] & x[22] & ~x[61] & ~x[63];
			partial_clause[336] 	= partial_clause_prev[336] & ~x[45];
			partial_clause[337] 	= partial_clause_prev[337] & ~x[10] & ~x[13] & ~x[36] & ~x[63];
			partial_clause[338] 	= partial_clause_prev[338] & 1'b1;
			partial_clause[339] 	= partial_clause_prev[339] & ~x[2] & ~x[11] & ~x[13] & ~x[32] & ~x[33] & ~x[35] & ~x[36] & ~x[42] & ~x[58];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[4] & ~x[9] & ~x[59] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[341] 	= partial_clause_prev[341] & 1'b1;
			partial_clause[342] 	= partial_clause_prev[342] & ~x[13] & ~x[29] & ~x[31] & ~x[37] & ~x[38] & ~x[39] & ~x[62];
			partial_clause[343] 	= partial_clause_prev[343] & ~x[7] & ~x[11] & ~x[15];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[10] & ~x[59] & ~x[61];
			partial_clause[345] 	= partial_clause_prev[345] & ~x[31] & ~x[61];
			partial_clause[346] 	= partial_clause_prev[346] & ~x[18] & ~x[19] & ~x[20] & ~x[32] & ~x[38] & ~x[39] & ~x[40] & ~x[41] & ~x[43] & ~x[44];
			partial_clause[347] 	= partial_clause_prev[347] & ~x[3] & ~x[10] & ~x[14] & ~x[15] & ~x[39] & ~x[44] & ~x[45];
			partial_clause[348] 	= partial_clause_prev[348] & ~x[33];
			partial_clause[349] 	= partial_clause_prev[349] & ~x[12];
			partial_clause[350] 	= partial_clause_prev[350] & ~x[1] & ~x[2] & ~x[3] & ~x[8] & ~x[10] & ~x[11] & ~x[12] & ~x[28] & ~x[29] & ~x[30] & ~x[31] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[38] & ~x[39] & ~x[41] & ~x[57] & ~x[58] & ~x[59] & ~x[60] & ~x[62];
			partial_clause[351] 	= partial_clause_prev[351] & 1'b1;
			partial_clause[352] 	= partial_clause_prev[352] & 1'b1;
			partial_clause[353] 	= partial_clause_prev[353] & ~x[48] & ~x[49];
			partial_clause[354] 	= partial_clause_prev[354] & ~x[3] & ~x[7] & ~x[61];
			partial_clause[355] 	= partial_clause_prev[355] & ~x[4] & ~x[7] & ~x[11] & ~x[38] & x[53];
			partial_clause[356] 	= partial_clause_prev[356] & ~x[7] & ~x[9] & ~x[35] & ~x[38] & ~x[39] & ~x[42] & ~x[44];
			partial_clause[357] 	= partial_clause_prev[357] & 1'b1;
			partial_clause[358] 	= partial_clause_prev[358] & ~x[11] & ~x[29] & ~x[36] & x[51] & ~x[58] & ~x[62];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[3] & ~x[33] & x[50] & x[51] & ~x[62];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[6] & ~x[9] & ~x[33] & ~x[34] & ~x[36] & ~x[38] & ~x[63];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[6] & ~x[7] & x[25] & ~x[33] & ~x[35] & ~x[57];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[10] & ~x[30] & ~x[32] & ~x[34];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[0] & ~x[8] & ~x[11] & ~x[13] & ~x[36] & ~x[37] & ~x[38] & ~x[43] & ~x[59] & ~x[60];
			partial_clause[364] 	= partial_clause_prev[364] & ~x[12];
			partial_clause[365] 	= partial_clause_prev[365] & 1'b1;
			partial_clause[366] 	= partial_clause_prev[366] & ~x[4] & ~x[7] & x[25] & ~x[33];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[5] & ~x[39];
			partial_clause[368] 	= partial_clause_prev[368] & 1'b1;
			partial_clause[369] 	= partial_clause_prev[369] & ~x[9] & ~x[32] & ~x[34] & ~x[35] & ~x[39] & ~x[61];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[2] & ~x[6] & ~x[7] & ~x[8] & ~x[15] & ~x[42] & ~x[63];
			partial_clause[371] 	= partial_clause_prev[371] & ~x[62];
			partial_clause[372] 	= partial_clause_prev[372] & ~x[9];
			partial_clause[373] 	= partial_clause_prev[373] & 1'b1;
			partial_clause[374] 	= partial_clause_prev[374] & ~x[63];
			partial_clause[375] 	= partial_clause_prev[375] & x[22];
			partial_clause[376] 	= partial_clause_prev[376] & ~x[1] & ~x[33] & ~x[40] & ~x[61];
			partial_clause[377] 	= partial_clause_prev[377] & ~x[6] & ~x[46];
			partial_clause[378] 	= partial_clause_prev[378] & ~x[1] & ~x[6] & ~x[9] & ~x[16] & ~x[63];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[5] & ~x[7] & ~x[13] & ~x[14];
			partial_clause[380] 	= partial_clause_prev[380] & ~x[3];
			partial_clause[381] 	= partial_clause_prev[381] & ~x[5] & ~x[7] & ~x[12] & ~x[36] & ~x[40] & ~x[41] & ~x[63];
			partial_clause[382] 	= partial_clause_prev[382] & 1'b1;
			partial_clause[383] 	= partial_clause_prev[383] & ~x[15] & ~x[36] & ~x[54] & ~x[55];
			partial_clause[384] 	= partial_clause_prev[384] & 1'b1;
			partial_clause[385] 	= partial_clause_prev[385] & ~x[41];
			partial_clause[386] 	= partial_clause_prev[386] & ~x[12] & ~x[22];
			partial_clause[387] 	= partial_clause_prev[387] & ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[17] & x[21] & ~x[27] & ~x[29] & ~x[35] & ~x[40] & ~x[56] & ~x[57] & ~x[58] & ~x[62] & ~x[63];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[9] & x[25] & ~x[36] & ~x[37];
			partial_clause[389] 	= partial_clause_prev[389] & 1'b1;
			partial_clause[390] 	= partial_clause_prev[390] & ~x[3] & ~x[7] & ~x[33] & ~x[58];
			partial_clause[391] 	= partial_clause_prev[391] & 1'b1;
			partial_clause[392] 	= partial_clause_prev[392] & x[22];
			partial_clause[393] 	= partial_clause_prev[393] & ~x[40];
			partial_clause[394] 	= partial_clause_prev[394] & ~x[4];
			partial_clause[395] 	= partial_clause_prev[395] & ~x[10] & ~x[38];
			partial_clause[396] 	= partial_clause_prev[396] & 1'b1;
			partial_clause[397] 	= partial_clause_prev[397] & ~x[1] & ~x[3];
			partial_clause[398] 	= partial_clause_prev[398] & 1'b1;
			partial_clause[399] 	= partial_clause_prev[399] & 1'b1;
			partial_clause[400] 	= partial_clause_prev[400] & ~x[1] & ~x[10] & ~x[40] & x[47] & ~x[57];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[1] & ~x[10] & ~x[11] & ~x[31] & ~x[34] & ~x[35] & ~x[42] & ~x[63];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[3] & ~x[12] & ~x[26] & ~x[38] & ~x[41];
			partial_clause[403] 	= partial_clause_prev[403] & ~x[11] & x[50];
			partial_clause[404] 	= partial_clause_prev[404] & 1'b1;
			partial_clause[405] 	= partial_clause_prev[405] & ~x[3] & ~x[4] & ~x[12] & ~x[13] & ~x[31] & ~x[35] & x[49];
			partial_clause[406] 	= partial_clause_prev[406] & ~x[5] & ~x[11] & ~x[12];
			partial_clause[407] 	= partial_clause_prev[407] & x[19] & ~x[61];
			partial_clause[408] 	= partial_clause_prev[408] & ~x[60];
			partial_clause[409] 	= partial_clause_prev[409] & ~x[1] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[8] & ~x[11] & ~x[13] & ~x[14] & ~x[32] & ~x[35] & ~x[38] & ~x[39] & ~x[58] & ~x[61];
			partial_clause[410] 	= partial_clause_prev[410] & ~x[4] & ~x[10] & ~x[33] & ~x[63];
			partial_clause[411] 	= partial_clause_prev[411] & ~x[4] & ~x[37];
			partial_clause[412] 	= partial_clause_prev[412] & ~x[2] & ~x[4] & ~x[8] & ~x[27] & ~x[30] & ~x[33] & ~x[37] & ~x[41] & ~x[55] & ~x[56] & ~x[60];
			partial_clause[413] 	= partial_clause_prev[413] & ~x[8] & ~x[14] & ~x[35];
			partial_clause[414] 	= partial_clause_prev[414] & ~x[4] & ~x[5] & ~x[6] & ~x[8] & ~x[11] & ~x[34];
			partial_clause[415] 	= partial_clause_prev[415] & 1'b1;
			partial_clause[416] 	= partial_clause_prev[416] & ~x[5] & ~x[12] & ~x[13] & ~x[36] & ~x[37] & ~x[58] & ~x[59] & ~x[61];
			partial_clause[417] 	= partial_clause_prev[417] & ~x[8];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[2] & ~x[6] & ~x[8] & ~x[11] & ~x[31] & ~x[32] & ~x[34] & ~x[38] & ~x[42] & ~x[43] & ~x[58] & ~x[60] & ~x[61];
			partial_clause[419] 	= partial_clause_prev[419] & x[21] & ~x[33];
			partial_clause[420] 	= partial_clause_prev[420] & ~x[17];
			partial_clause[421] 	= partial_clause_prev[421] & ~x[3] & ~x[5] & ~x[12] & ~x[38];
			partial_clause[422] 	= partial_clause_prev[422] & ~x[8] & ~x[12] & ~x[14] & ~x[17] & ~x[18] & ~x[62] & ~x[63];
			partial_clause[423] 	= partial_clause_prev[423] & ~x[33] & ~x[37];
			partial_clause[424] 	= partial_clause_prev[424] & ~x[7] & ~x[40];
			partial_clause[425] 	= partial_clause_prev[425] & ~x[20] & ~x[24] & ~x[49] & ~x[51];
			partial_clause[426] 	= partial_clause_prev[426] & ~x[2] & ~x[6] & ~x[7] & ~x[10] & ~x[36] & ~x[39] & ~x[41] & ~x[55] & ~x[56];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[0] & ~x[6] & ~x[7] & ~x[38] & ~x[57] & ~x[62];
			partial_clause[428] 	= partial_clause_prev[428] & 1'b1;
			partial_clause[429] 	= partial_clause_prev[429] & 1'b1;
			partial_clause[430] 	= partial_clause_prev[430] & ~x[4] & ~x[7] & ~x[13] & ~x[15] & ~x[17] & ~x[30] & ~x[32] & ~x[39] & ~x[44] & ~x[60] & ~x[63];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[3] & ~x[34] & ~x[38];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[1] & ~x[4] & ~x[8] & ~x[15] & ~x[36] & ~x[60];
			partial_clause[433] 	= partial_clause_prev[433] & ~x[19] & ~x[48] & ~x[62];
			partial_clause[434] 	= partial_clause_prev[434] & x[26] & x[54] & ~x[61];
			partial_clause[435] 	= partial_clause_prev[435] & ~x[4] & ~x[7] & ~x[11] & ~x[16] & ~x[32] & ~x[35] & ~x[37] & ~x[40] & ~x[41] & ~x[42] & ~x[58] & ~x[60] & ~x[61] & ~x[63];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[4] & ~x[6] & ~x[7] & ~x[10] & ~x[33] & ~x[36];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[7] & ~x[8] & ~x[33] & ~x[36] & ~x[37] & ~x[39] & ~x[62];
			partial_clause[438] 	= partial_clause_prev[438] & ~x[1] & x[24];
			partial_clause[439] 	= partial_clause_prev[439] & ~x[37];
			partial_clause[440] 	= partial_clause_prev[440] & ~x[42];
			partial_clause[441] 	= partial_clause_prev[441] & ~x[39] & ~x[41] & ~x[42];
			partial_clause[442] 	= partial_clause_prev[442] & ~x[20] & ~x[47];
			partial_clause[443] 	= partial_clause_prev[443] & ~x[2] & ~x[4] & ~x[10] & ~x[28] & ~x[29] & ~x[31] & ~x[36] & ~x[39] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[444] 	= partial_clause_prev[444] & ~x[50];
			partial_clause[445] 	= partial_clause_prev[445] & ~x[12] & ~x[19] & ~x[46];
			partial_clause[446] 	= partial_clause_prev[446] & ~x[6] & ~x[8] & ~x[11] & ~x[31] & ~x[35] & ~x[40] & ~x[62];
			partial_clause[447] 	= partial_clause_prev[447] & ~x[2] & ~x[9] & ~x[14] & ~x[31] & ~x[36] & ~x[61];
			partial_clause[448] 	= partial_clause_prev[448] & ~x[20] & ~x[48];
			partial_clause[449] 	= partial_clause_prev[449] & ~x[13] & ~x[30] & ~x[36] & ~x[59] & ~x[63];
			partial_clause[450] 	= partial_clause_prev[450] & ~x[8] & ~x[9] & ~x[35] & ~x[38];
			partial_clause[451] 	= partial_clause_prev[451] & ~x[55];
			partial_clause[452] 	= partial_clause_prev[452] & ~x[13] & x[24] & ~x[27];
			partial_clause[453] 	= partial_clause_prev[453] & ~x[59] & ~x[61];
			partial_clause[454] 	= partial_clause_prev[454] & ~x[7] & ~x[33] & ~x[39] & ~x[61];
			partial_clause[455] 	= partial_clause_prev[455] & ~x[5] & ~x[8] & ~x[9] & ~x[10] & x[24] & ~x[37] & ~x[38];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[7] & ~x[13] & ~x[14] & ~x[29] & ~x[34] & ~x[36] & ~x[44] & ~x[60];
			partial_clause[457] 	= partial_clause_prev[457] & ~x[36];
			partial_clause[458] 	= partial_clause_prev[458] & ~x[13] & ~x[14] & ~x[15] & ~x[34] & ~x[39];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[11] & ~x[62];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[5] & ~x[6] & ~x[9] & ~x[32] & ~x[35] & ~x[37] & ~x[40];
			partial_clause[461] 	= partial_clause_prev[461] & ~x[3] & ~x[29] & ~x[33];
			partial_clause[462] 	= partial_clause_prev[462] & ~x[0] & ~x[36];
			partial_clause[463] 	= partial_clause_prev[463] & ~x[13] & ~x[14] & ~x[16] & ~x[42];
			partial_clause[464] 	= partial_clause_prev[464] & ~x[5] & ~x[30] & ~x[32];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[3] & ~x[5] & ~x[6] & ~x[18] & x[22] & ~x[31] & x[50] & ~x[55] & ~x[59];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[5] & ~x[7] & ~x[11] & ~x[12] & ~x[34] & ~x[35] & ~x[50] & ~x[51];
			partial_clause[467] 	= partial_clause_prev[467] & ~x[0] & ~x[18] & ~x[19] & ~x[42];
			partial_clause[468] 	= partial_clause_prev[468] & ~x[4] & ~x[38] & ~x[40] & ~x[59] & ~x[61] & ~x[62];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[2] & ~x[5] & ~x[12] & ~x[18] & ~x[39] & ~x[45] & ~x[46];
			partial_clause[470] 	= partial_clause_prev[470] & ~x[15] & x[50];
			partial_clause[471] 	= partial_clause_prev[471] & ~x[10] & ~x[11] & ~x[15] & ~x[41] & ~x[59];
			partial_clause[472] 	= partial_clause_prev[472] & ~x[31] & ~x[35];
			partial_clause[473] 	= partial_clause_prev[473] & ~x[5] & ~x[6] & ~x[10] & ~x[13] & ~x[37] & ~x[38];
			partial_clause[474] 	= partial_clause_prev[474] & ~x[15] & ~x[43];
			partial_clause[475] 	= partial_clause_prev[475] & ~x[5] & ~x[11] & ~x[31] & ~x[40] & ~x[56] & ~x[58] & ~x[61];
			partial_clause[476] 	= partial_clause_prev[476] & ~x[10];
			partial_clause[477] 	= partial_clause_prev[477] & ~x[37] & ~x[38] & ~x[39];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[6] & ~x[32];
			partial_clause[479] 	= partial_clause_prev[479] & 1'b1;
			partial_clause[480] 	= partial_clause_prev[480] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[16] & ~x[17] & ~x[18] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[38] & ~x[39] & ~x[40] & ~x[43] & ~x[44] & ~x[45] & ~x[57] & ~x[58] & ~x[59] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[481] 	= partial_clause_prev[481] & 1'b1;
			partial_clause[482] 	= partial_clause_prev[482] & ~x[17] & ~x[39] & ~x[42];
			partial_clause[483] 	= partial_clause_prev[483] & ~x[57];
			partial_clause[484] 	= partial_clause_prev[484] & ~x[42];
			partial_clause[485] 	= partial_clause_prev[485] & x[57];
			partial_clause[486] 	= partial_clause_prev[486] & ~x[7] & ~x[34];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[8] & ~x[34] & ~x[38] & ~x[62];
			partial_clause[488] 	= partial_clause_prev[488] & ~x[39];
			partial_clause[489] 	= partial_clause_prev[489] & 1'b1;
			partial_clause[490] 	= partial_clause_prev[490] & ~x[25];
			partial_clause[491] 	= partial_clause_prev[491] & ~x[6] & x[51];
			partial_clause[492] 	= partial_clause_prev[492] & ~x[2] & ~x[3] & ~x[10] & ~x[37];
			partial_clause[493] 	= partial_clause_prev[493] & x[51];
			partial_clause[494] 	= partial_clause_prev[494] & 1'b1;
			partial_clause[495] 	= partial_clause_prev[495] & ~x[9] & ~x[10] & ~x[60];
			partial_clause[496] 	= partial_clause_prev[496] & 1'b1;
			partial_clause[497] 	= partial_clause_prev[497] & ~x[48];
			partial_clause[498] 	= partial_clause_prev[498] & 1'b1;
			partial_clause[499] 	= partial_clause_prev[499] & 1'b1;
		end
	end
endmodule


module HCB_7 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[4] & ~x[24] & ~x[51] & ~x[53] & ~x[55] & ~x[58] & ~x[59];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[3] & ~x[4] & ~x[26] & ~x[27] & ~x[33] & ~x[53] & ~x[62];
			partial_clause[2] 	= partial_clause_prev[2] & ~x[32] & ~x[33] & ~x[35] & ~x[37] & ~x[52] & ~x[54];
			partial_clause[3] 	= partial_clause_prev[3] & ~x[4] & ~x[23] & ~x[49] & ~x[53];
			partial_clause[4] 	= partial_clause_prev[4] & ~x[29] & ~x[30] & ~x[53];
			partial_clause[5] 	= partial_clause_prev[5] & ~x[1] & ~x[23] & ~x[30] & ~x[54] & ~x[59] & ~x[61];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[4] & ~x[25] & ~x[26] & ~x[27] & ~x[53] & ~x[54];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[5] & ~x[54];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[26] & ~x[29];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[3] & ~x[7] & ~x[8] & ~x[28] & ~x[31] & ~x[32] & ~x[35] & ~x[36] & ~x[37] & ~x[50] & ~x[52] & ~x[60];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[5] & ~x[6] & ~x[24] & ~x[28] & ~x[32] & ~x[61];
			partial_clause[11] 	= partial_clause_prev[11] & ~x[3] & ~x[23] & ~x[24] & ~x[25] & ~x[26] & ~x[30] & ~x[55];
			partial_clause[12] 	= partial_clause_prev[12] & x[16] & ~x[25] & ~x[30] & ~x[55] & ~x[59];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[2] & ~x[3] & ~x[47] & ~x[49] & ~x[50] & ~x[56] & ~x[58];
			partial_clause[14] 	= partial_clause_prev[14] & ~x[39];
			partial_clause[15] 	= partial_clause_prev[15] & 1'b1;
			partial_clause[16] 	= partial_clause_prev[16] & ~x[1] & ~x[57];
			partial_clause[17] 	= partial_clause_prev[17] & 1'b1;
			partial_clause[18] 	= partial_clause_prev[18] & x[11];
			partial_clause[19] 	= partial_clause_prev[19] & ~x[0] & ~x[25] & ~x[37] & ~x[38] & ~x[40] & ~x[56];
			partial_clause[20] 	= partial_clause_prev[20] & x[18] & ~x[26] & x[46] & ~x[56];
			partial_clause[21] 	= partial_clause_prev[21] & ~x[6] & ~x[8] & ~x[54];
			partial_clause[22] 	= partial_clause_prev[22] & ~x[27] & ~x[28];
			partial_clause[23] 	= partial_clause_prev[23] & ~x[1] & ~x[4] & ~x[27] & ~x[28] & ~x[31] & ~x[55] & ~x[56];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[0] & ~x[2] & ~x[3] & ~x[4] & ~x[16] & ~x[17] & ~x[25] & ~x[27] & ~x[32] & ~x[53] & ~x[54] & ~x[56] & ~x[58] & ~x[59] & ~x[61];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[0] & ~x[1] & ~x[2] & ~x[6] & ~x[27] & ~x[29] & ~x[32] & ~x[34] & ~x[49] & ~x[53] & ~x[55] & ~x[56];
			partial_clause[26] 	= partial_clause_prev[26] & 1'b1;
			partial_clause[27] 	= partial_clause_prev[27] & ~x[1] & ~x[3] & ~x[25] & ~x[54];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[2] & ~x[4] & ~x[46] & ~x[57] & ~x[60];
			partial_clause[29] 	= partial_clause_prev[29] & ~x[3] & ~x[4] & ~x[26];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[0] & ~x[25] & ~x[30];
			partial_clause[31] 	= partial_clause_prev[31] & ~x[26] & ~x[30] & ~x[31] & ~x[33] & ~x[54] & ~x[58];
			partial_clause[32] 	= partial_clause_prev[32] & 1'b1;
			partial_clause[33] 	= partial_clause_prev[33] & ~x[17];
			partial_clause[34] 	= partial_clause_prev[34] & ~x[28] & ~x[29] & ~x[30] & ~x[54] & ~x[57] & ~x[59];
			partial_clause[35] 	= partial_clause_prev[35] & ~x[12] & ~x[15] & ~x[26] & ~x[30] & ~x[39] & ~x[42];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[1] & ~x[4] & ~x[9] & ~x[21] & ~x[49] & ~x[52] & ~x[60];
			partial_clause[37] 	= partial_clause_prev[37] & ~x[5];
			partial_clause[38] 	= partial_clause_prev[38] & ~x[0] & ~x[1] & ~x[27] & ~x[58];
			partial_clause[39] 	= partial_clause_prev[39] & ~x[21] & ~x[32] & ~x[45] & ~x[46] & ~x[49];
			partial_clause[40] 	= partial_clause_prev[40] & ~x[28] & ~x[53];
			partial_clause[41] 	= partial_clause_prev[41] & x[38];
			partial_clause[42] 	= partial_clause_prev[42] & 1'b1;
			partial_clause[43] 	= partial_clause_prev[43] & ~x[5] & x[13] & ~x[29] & ~x[33];
			partial_clause[44] 	= partial_clause_prev[44] & ~x[15] & ~x[45] & ~x[46];
			partial_clause[45] 	= partial_clause_prev[45] & ~x[30] & ~x[31] & ~x[46] & ~x[47] & ~x[58] & ~x[59] & ~x[60];
			partial_clause[46] 	= partial_clause_prev[46] & ~x[0] & ~x[6] & ~x[22] & ~x[24] & ~x[31] & ~x[53] & ~x[54] & ~x[56];
			partial_clause[47] 	= partial_clause_prev[47] & ~x[26] & ~x[50] & ~x[59] & ~x[60] & ~x[62];
			partial_clause[48] 	= partial_clause_prev[48] & 1'b1;
			partial_clause[49] 	= partial_clause_prev[49] & ~x[61];
			partial_clause[50] 	= partial_clause_prev[50] & ~x[27];
			partial_clause[51] 	= partial_clause_prev[51] & 1'b1;
			partial_clause[52] 	= partial_clause_prev[52] & 1'b1;
			partial_clause[53] 	= partial_clause_prev[53] & ~x[20];
			partial_clause[54] 	= partial_clause_prev[54] & 1'b1;
			partial_clause[55] 	= partial_clause_prev[55] & x[38];
			partial_clause[56] 	= partial_clause_prev[56] & 1'b1;
			partial_clause[57] 	= partial_clause_prev[57] & ~x[4] & ~x[32] & ~x[55] & ~x[58];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[4] & ~x[6] & ~x[22] & ~x[23] & ~x[26] & ~x[29] & ~x[31] & ~x[34] & ~x[51] & ~x[57];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[0] & ~x[25] & ~x[26] & ~x[53] & ~x[54] & ~x[55] & ~x[57];
			partial_clause[60] 	= partial_clause_prev[60] & ~x[33] & ~x[36] & ~x[62];
			partial_clause[61] 	= partial_clause_prev[61] & ~x[44];
			partial_clause[62] 	= partial_clause_prev[62] & ~x[0] & ~x[29] & ~x[33] & ~x[38] & ~x[39] & ~x[50] & ~x[52];
			partial_clause[63] 	= partial_clause_prev[63] & ~x[3] & ~x[28] & ~x[32] & ~x[59];
			partial_clause[64] 	= partial_clause_prev[64] & 1'b1;
			partial_clause[65] 	= partial_clause_prev[65] & 1'b1;
			partial_clause[66] 	= partial_clause_prev[66] & 1'b1;
			partial_clause[67] 	= partial_clause_prev[67] & 1'b1;
			partial_clause[68] 	= partial_clause_prev[68] & ~x[11] & ~x[14] & ~x[27] & ~x[56];
			partial_clause[69] 	= partial_clause_prev[69] & ~x[7] & ~x[21] & ~x[35] & ~x[37] & ~x[52] & ~x[53];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[3] & ~x[20] & ~x[21] & ~x[31] & ~x[45];
			partial_clause[71] 	= partial_clause_prev[71] & ~x[6] & ~x[31] & ~x[36];
			partial_clause[72] 	= partial_clause_prev[72] & 1'b1;
			partial_clause[73] 	= partial_clause_prev[73] & 1'b1;
			partial_clause[74] 	= partial_clause_prev[74] & ~x[9] & ~x[10] & ~x[39] & ~x[40];
			partial_clause[75] 	= partial_clause_prev[75] & ~x[34] & ~x[36] & ~x[52] & ~x[62];
			partial_clause[76] 	= partial_clause_prev[76] & ~x[1] & ~x[3] & ~x[28] & ~x[33] & ~x[49] & ~x[58] & ~x[59];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[5];
			partial_clause[78] 	= partial_clause_prev[78] & ~x[34];
			partial_clause[79] 	= partial_clause_prev[79] & ~x[30] & ~x[59] & ~x[61];
			partial_clause[80] 	= partial_clause_prev[80] & ~x[26];
			partial_clause[81] 	= partial_clause_prev[81] & x[13] & ~x[20];
			partial_clause[82] 	= partial_clause_prev[82] & x[8] & ~x[58];
			partial_clause[83] 	= partial_clause_prev[83] & 1'b1;
			partial_clause[84] 	= partial_clause_prev[84] & ~x[22] & ~x[27] & ~x[35] & ~x[60];
			partial_clause[85] 	= partial_clause_prev[85] & ~x[1] & ~x[4] & ~x[22] & ~x[26] & ~x[29] & ~x[32] & ~x[53];
			partial_clause[86] 	= partial_clause_prev[86] & ~x[0] & ~x[30];
			partial_clause[87] 	= partial_clause_prev[87] & ~x[27];
			partial_clause[88] 	= partial_clause_prev[88] & ~x[26] & ~x[28] & ~x[41] & ~x[42] & ~x[55] & ~x[58] & ~x[59];
			partial_clause[89] 	= partial_clause_prev[89] & ~x[1] & ~x[5] & ~x[9] & ~x[53] & ~x[63];
			partial_clause[90] 	= partial_clause_prev[90] & 1'b1;
			partial_clause[91] 	= partial_clause_prev[91] & ~x[33] & ~x[35];
			partial_clause[92] 	= partial_clause_prev[92] & ~x[0] & ~x[4] & ~x[27] & ~x[50];
			partial_clause[93] 	= partial_clause_prev[93] & ~x[0] & ~x[1] & ~x[2] & ~x[4] & ~x[5] & ~x[23] & ~x[26] & ~x[27] & ~x[29] & ~x[30] & ~x[31] & ~x[32] & ~x[34] & ~x[35] & ~x[60] & ~x[61];
			partial_clause[94] 	= partial_clause_prev[94] & ~x[13] & ~x[40];
			partial_clause[95] 	= partial_clause_prev[95] & ~x[1] & ~x[8] & ~x[19] & ~x[20] & ~x[22] & ~x[23] & ~x[29] & ~x[52] & ~x[53] & ~x[56] & ~x[57] & ~x[61] & ~x[62];
			partial_clause[96] 	= partial_clause_prev[96] & ~x[12] & ~x[39];
			partial_clause[97] 	= partial_clause_prev[97] & ~x[1] & ~x[2] & ~x[4] & ~x[6] & ~x[7] & ~x[21] & ~x[22] & ~x[25] & ~x[29] & ~x[33] & ~x[50] & ~x[52] & ~x[54] & ~x[58] & ~x[59] & ~x[61];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[2] & ~x[27] & ~x[30] & ~x[55] & ~x[57];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[1] & ~x[2] & ~x[3] & ~x[5] & ~x[6] & ~x[23] & ~x[25] & ~x[27] & ~x[30] & ~x[34] & ~x[52] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[59] & ~x[60] & ~x[62];
			partial_clause[100] 	= partial_clause_prev[100] & x[11] & x[38];
			partial_clause[101] 	= partial_clause_prev[101] & 1'b1;
			partial_clause[102] 	= partial_clause_prev[102] & ~x[18] & ~x[19];
			partial_clause[103] 	= partial_clause_prev[103] & ~x[0] & ~x[21] & ~x[23] & ~x[24] & ~x[26] & ~x[30] & ~x[54] & ~x[56] & ~x[58];
			partial_clause[104] 	= partial_clause_prev[104] & ~x[27] & ~x[60];
			partial_clause[105] 	= partial_clause_prev[105] & ~x[1] & ~x[53] & ~x[57] & ~x[59] & ~x[60];
			partial_clause[106] 	= partial_clause_prev[106] & ~x[25] & ~x[26] & ~x[31] & ~x[56] & ~x[59];
			partial_clause[107] 	= partial_clause_prev[107] & ~x[2] & ~x[27] & ~x[29] & ~x[58] & ~x[60] & ~x[61];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[2] & ~x[4] & x[16] & ~x[28] & ~x[31] & ~x[57] & ~x[60] & ~x[61];
			partial_clause[109] 	= partial_clause_prev[109] & 1'b1;
			partial_clause[110] 	= partial_clause_prev[110] & x[42];
			partial_clause[111] 	= partial_clause_prev[111] & 1'b1;
			partial_clause[112] 	= partial_clause_prev[112] & ~x[25] & ~x[26] & ~x[33] & ~x[39] & ~x[40];
			partial_clause[113] 	= partial_clause_prev[113] & ~x[2];
			partial_clause[114] 	= partial_clause_prev[114] & 1'b1;
			partial_clause[115] 	= partial_clause_prev[115] & ~x[2] & ~x[4] & ~x[5] & ~x[23] & ~x[27] & ~x[51] & ~x[57];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[1] & ~x[5] & ~x[25] & ~x[48] & ~x[62];
			partial_clause[117] 	= partial_clause_prev[117] & 1'b1;
			partial_clause[118] 	= partial_clause_prev[118] & ~x[5] & ~x[10] & ~x[22] & ~x[29] & ~x[32] & ~x[35] & ~x[52];
			partial_clause[119] 	= partial_clause_prev[119] & ~x[1] & ~x[25] & ~x[27] & ~x[29] & ~x[32] & ~x[34] & ~x[49] & ~x[56] & ~x[59] & ~x[61] & ~x[62];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[4] & ~x[24] & ~x[25] & ~x[26] & ~x[31] & ~x[32] & ~x[33] & ~x[53] & ~x[54] & ~x[58] & ~x[59] & ~x[60];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[0];
			partial_clause[122] 	= partial_clause_prev[122] & ~x[18] & ~x[31] & ~x[48];
			partial_clause[123] 	= partial_clause_prev[123] & ~x[2] & ~x[25] & ~x[28] & ~x[53] & ~x[56] & ~x[58];
			partial_clause[124] 	= partial_clause_prev[124] & ~x[16] & x[47] & ~x[53];
			partial_clause[125] 	= partial_clause_prev[125] & x[40];
			partial_clause[126] 	= partial_clause_prev[126] & ~x[1] & ~x[3] & ~x[62];
			partial_clause[127] 	= partial_clause_prev[127] & ~x[2] & ~x[4] & ~x[5] & ~x[6] & x[15] & ~x[20] & ~x[21] & ~x[28] & ~x[29] & ~x[30] & ~x[32] & ~x[35] & ~x[51] & ~x[55] & ~x[56] & ~x[60];
			partial_clause[128] 	= partial_clause_prev[128] & ~x[2] & ~x[26];
			partial_clause[129] 	= partial_clause_prev[129] & ~x[1] & ~x[4] & ~x[26] & ~x[28] & ~x[32];
			partial_clause[130] 	= partial_clause_prev[130] & ~x[28];
			partial_clause[131] 	= partial_clause_prev[131] & ~x[34];
			partial_clause[132] 	= partial_clause_prev[132] & ~x[0] & ~x[4] & ~x[27];
			partial_clause[133] 	= partial_clause_prev[133] & x[42];
			partial_clause[134] 	= partial_clause_prev[134] & ~x[1] & ~x[4] & ~x[5] & ~x[21] & ~x[24] & ~x[25] & ~x[28] & ~x[29] & ~x[30] & ~x[31] & ~x[34] & ~x[38] & ~x[52] & ~x[58];
			partial_clause[135] 	= partial_clause_prev[135] & ~x[1] & ~x[52] & ~x[55];
			partial_clause[136] 	= partial_clause_prev[136] & ~x[8] & ~x[28] & ~x[35] & ~x[37] & ~x[39] & ~x[40] & ~x[41] & ~x[51] & ~x[54] & ~x[56] & ~x[57];
			partial_clause[137] 	= partial_clause_prev[137] & 1'b1;
			partial_clause[138] 	= partial_clause_prev[138] & ~x[35];
			partial_clause[139] 	= partial_clause_prev[139] & ~x[2] & ~x[3] & ~x[25] & ~x[29] & ~x[30] & ~x[31] & ~x[33] & ~x[53] & ~x[56] & ~x[57] & ~x[61];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[21] & ~x[22] & ~x[26] & ~x[29] & ~x[31] & ~x[33] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[60] & ~x[62];
			partial_clause[141] 	= partial_clause_prev[141] & ~x[51] & ~x[59] & ~x[62];
			partial_clause[142] 	= partial_clause_prev[142] & ~x[0] & ~x[3] & ~x[5] & ~x[8] & ~x[20] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & ~x[30] & ~x[50] & ~x[52] & ~x[56] & ~x[61];
			partial_clause[143] 	= partial_clause_prev[143] & 1'b1;
			partial_clause[144] 	= partial_clause_prev[144] & ~x[29];
			partial_clause[145] 	= partial_clause_prev[145] & 1'b1;
			partial_clause[146] 	= partial_clause_prev[146] & ~x[0] & ~x[3] & ~x[17] & ~x[18] & ~x[25] & ~x[30] & ~x[31] & ~x[46] & ~x[47];
			partial_clause[147] 	= partial_clause_prev[147] & ~x[1] & ~x[2] & ~x[25] & ~x[27] & ~x[28];
			partial_clause[148] 	= partial_clause_prev[148] & x[15] & ~x[28] & x[43] & ~x[62];
			partial_clause[149] 	= partial_clause_prev[149] & 1'b1;
			partial_clause[150] 	= partial_clause_prev[150] & ~x[0] & ~x[23] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[59];
			partial_clause[151] 	= partial_clause_prev[151] & 1'b1;
			partial_clause[152] 	= partial_clause_prev[152] & x[19] & ~x[25] & x[45] & ~x[53];
			partial_clause[153] 	= partial_clause_prev[153] & ~x[1] & ~x[28] & ~x[32] & ~x[33] & ~x[43] & ~x[54] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[154] 	= partial_clause_prev[154] & ~x[9] & x[13] & ~x[52];
			partial_clause[155] 	= partial_clause_prev[155] & 1'b1;
			partial_clause[156] 	= partial_clause_prev[156] & 1'b1;
			partial_clause[157] 	= partial_clause_prev[157] & 1'b1;
			partial_clause[158] 	= partial_clause_prev[158] & ~x[3] & ~x[4] & ~x[19] & ~x[20] & ~x[21] & ~x[26] & ~x[28] & ~x[29] & ~x[30] & ~x[46] & ~x[47] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[54] & ~x[55] & ~x[59];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[3] & ~x[6] & ~x[18] & ~x[29] & ~x[34] & ~x[58] & ~x[60] & ~x[61];
			partial_clause[160] 	= partial_clause_prev[160] & ~x[8] & ~x[56];
			partial_clause[161] 	= partial_clause_prev[161] & ~x[4] & ~x[23] & ~x[28] & ~x[29];
			partial_clause[162] 	= partial_clause_prev[162] & ~x[0] & ~x[3] & ~x[53] & ~x[54] & ~x[58];
			partial_clause[163] 	= partial_clause_prev[163] & 1'b1;
			partial_clause[164] 	= partial_clause_prev[164] & ~x[30] & ~x[39];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[27] & ~x[29] & ~x[51] & ~x[54] & ~x[55] & ~x[56] & ~x[59] & ~x[62] & ~x[63];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[19] & ~x[25] & ~x[26];
			partial_clause[167] 	= partial_clause_prev[167] & 1'b1;
			partial_clause[168] 	= partial_clause_prev[168] & ~x[3] & ~x[25] & ~x[58];
			partial_clause[169] 	= partial_clause_prev[169] & ~x[56];
			partial_clause[170] 	= partial_clause_prev[170] & ~x[25];
			partial_clause[171] 	= partial_clause_prev[171] & ~x[0] & ~x[2] & ~x[5] & ~x[21] & ~x[26] & ~x[27] & ~x[29] & ~x[32] & ~x[51];
			partial_clause[172] 	= partial_clause_prev[172] & 1'b1;
			partial_clause[173] 	= partial_clause_prev[173] & ~x[27] & ~x[53] & ~x[58];
			partial_clause[174] 	= partial_clause_prev[174] & ~x[0];
			partial_clause[175] 	= partial_clause_prev[175] & 1'b1;
			partial_clause[176] 	= partial_clause_prev[176] & 1'b1;
			partial_clause[177] 	= partial_clause_prev[177] & ~x[3] & ~x[23] & ~x[33] & ~x[51] & ~x[53];
			partial_clause[178] 	= partial_clause_prev[178] & ~x[2] & ~x[21] & ~x[48];
			partial_clause[179] 	= partial_clause_prev[179] & 1'b1;
			partial_clause[180] 	= partial_clause_prev[180] & ~x[34];
			partial_clause[181] 	= partial_clause_prev[181] & x[11];
			partial_clause[182] 	= partial_clause_prev[182] & x[45];
			partial_clause[183] 	= partial_clause_prev[183] & ~x[3] & ~x[4] & ~x[6] & ~x[7] & ~x[25] & ~x[28] & ~x[29] & ~x[37] & ~x[49] & ~x[54] & ~x[58];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[6] & ~x[20] & ~x[23] & ~x[25] & ~x[27] & ~x[29] & ~x[34] & ~x[57] & ~x[60] & ~x[61];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[1] & ~x[24] & ~x[52] & ~x[55];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[2] & ~x[4] & ~x[22] & ~x[32] & ~x[52] & ~x[56] & ~x[58] & ~x[60] & ~x[62];
			partial_clause[187] 	= partial_clause_prev[187] & ~x[2] & ~x[25] & ~x[50] & ~x[55];
			partial_clause[188] 	= partial_clause_prev[188] & ~x[44] & ~x[53];
			partial_clause[189] 	= partial_clause_prev[189] & ~x[12];
			partial_clause[190] 	= partial_clause_prev[190] & x[16] & ~x[20] & ~x[48] & ~x[51] & ~x[55];
			partial_clause[191] 	= partial_clause_prev[191] & ~x[24];
			partial_clause[192] 	= partial_clause_prev[192] & ~x[1] & ~x[58];
			partial_clause[193] 	= partial_clause_prev[193] & ~x[3] & ~x[5] & ~x[22] & ~x[23] & ~x[24] & ~x[32] & ~x[35] & ~x[57];
			partial_clause[194] 	= partial_clause_prev[194] & ~x[24] & ~x[32];
			partial_clause[195] 	= partial_clause_prev[195] & ~x[1] & ~x[2] & ~x[26] & ~x[27] & ~x[33] & ~x[47] & ~x[50] & ~x[54] & ~x[56];
			partial_clause[196] 	= partial_clause_prev[196] & 1'b1;
			partial_clause[197] 	= partial_clause_prev[197] & ~x[0] & ~x[26] & ~x[29] & ~x[31] & ~x[32] & ~x[34] & ~x[55];
			partial_clause[198] 	= partial_clause_prev[198] & 1'b1;
			partial_clause[199] 	= partial_clause_prev[199] & 1'b1;
			partial_clause[200] 	= partial_clause_prev[200] & ~x[31] & ~x[42];
			partial_clause[201] 	= partial_clause_prev[201] & ~x[27] & ~x[54] & ~x[55] & ~x[57] & ~x[58] & ~x[60];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[1] & ~x[4] & ~x[9] & ~x[27] & ~x[31] & ~x[55] & ~x[63];
			partial_clause[203] 	= partial_clause_prev[203] & ~x[51];
			partial_clause[204] 	= partial_clause_prev[204] & ~x[2] & ~x[21] & ~x[30] & ~x[48] & ~x[52] & ~x[57] & ~x[61];
			partial_clause[205] 	= partial_clause_prev[205] & 1'b1;
			partial_clause[206] 	= partial_clause_prev[206] & ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[28] & ~x[29] & ~x[31];
			partial_clause[207] 	= partial_clause_prev[207] & ~x[6] & ~x[29] & ~x[54] & ~x[58] & ~x[60] & ~x[62];
			partial_clause[208] 	= partial_clause_prev[208] & ~x[28] & ~x[52] & ~x[60];
			partial_clause[209] 	= partial_clause_prev[209] & 1'b1;
			partial_clause[210] 	= partial_clause_prev[210] & ~x[57];
			partial_clause[211] 	= partial_clause_prev[211] & ~x[38];
			partial_clause[212] 	= partial_clause_prev[212] & ~x[25] & ~x[29] & ~x[31] & ~x[53];
			partial_clause[213] 	= partial_clause_prev[213] & 1'b1;
			partial_clause[214] 	= partial_clause_prev[214] & x[10];
			partial_clause[215] 	= partial_clause_prev[215] & x[9];
			partial_clause[216] 	= partial_clause_prev[216] & ~x[56];
			partial_clause[217] 	= partial_clause_prev[217] & 1'b1;
			partial_clause[218] 	= partial_clause_prev[218] & ~x[19] & ~x[47];
			partial_clause[219] 	= partial_clause_prev[219] & ~x[4] & ~x[57];
			partial_clause[220] 	= partial_clause_prev[220] & ~x[3] & ~x[4] & ~x[20] & ~x[29] & ~x[32] & ~x[51] & ~x[58];
			partial_clause[221] 	= partial_clause_prev[221] & ~x[61];
			partial_clause[222] 	= partial_clause_prev[222] & 1'b1;
			partial_clause[223] 	= partial_clause_prev[223] & ~x[22] & ~x[31];
			partial_clause[224] 	= partial_clause_prev[224] & ~x[1] & ~x[29] & ~x[50] & ~x[54] & ~x[57] & ~x[58];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[58];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[25] & ~x[26] & ~x[27] & ~x[56] & ~x[57] & ~x[59];
			partial_clause[227] 	= partial_clause_prev[227] & ~x[29];
			partial_clause[228] 	= partial_clause_prev[228] & ~x[1] & ~x[3] & ~x[4] & ~x[26] & ~x[30] & ~x[32] & ~x[47] & ~x[58] & ~x[59];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[5] & ~x[24] & ~x[28] & ~x[52] & ~x[61];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[0] & ~x[1] & ~x[6] & ~x[24] & ~x[25] & ~x[27] & ~x[28] & ~x[30] & ~x[31] & ~x[33] & ~x[49] & ~x[51] & ~x[54] & ~x[57];
			partial_clause[231] 	= partial_clause_prev[231] & ~x[27] & ~x[29] & ~x[53];
			partial_clause[232] 	= partial_clause_prev[232] & 1'b1;
			partial_clause[233] 	= partial_clause_prev[233] & x[18] & ~x[23] & ~x[57];
			partial_clause[234] 	= partial_clause_prev[234] & ~x[2];
			partial_clause[235] 	= partial_clause_prev[235] & ~x[12] & ~x[13];
			partial_clause[236] 	= partial_clause_prev[236] & ~x[9] & ~x[20] & ~x[27] & ~x[37];
			partial_clause[237] 	= partial_clause_prev[237] & ~x[29];
			partial_clause[238] 	= partial_clause_prev[238] & x[15] & ~x[32] & ~x[37] & ~x[62];
			partial_clause[239] 	= partial_clause_prev[239] & x[41] & x[42] & ~x[47];
			partial_clause[240] 	= partial_clause_prev[240] & ~x[18] & ~x[21] & ~x[27] & x[43] & ~x[54] & ~x[58];
			partial_clause[241] 	= partial_clause_prev[241] & ~x[22] & ~x[23];
			partial_clause[242] 	= partial_clause_prev[242] & ~x[1] & ~x[3] & ~x[4] & ~x[25] & ~x[29] & ~x[31] & ~x[50] & ~x[51] & ~x[55];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[32] & ~x[59] & ~x[60];
			partial_clause[244] 	= partial_clause_prev[244] & ~x[60];
			partial_clause[245] 	= partial_clause_prev[245] & 1'b1;
			partial_clause[246] 	= partial_clause_prev[246] & ~x[30] & ~x[53] & ~x[55];
			partial_clause[247] 	= partial_clause_prev[247] & ~x[0] & ~x[2] & ~x[7] & ~x[22] & ~x[27] & ~x[31] & ~x[34] & ~x[48] & ~x[49] & ~x[56] & ~x[60];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[2] & ~x[4] & ~x[5] & ~x[23] & ~x[25] & ~x[26] & ~x[34] & ~x[56] & ~x[58] & ~x[60];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[39] & ~x[60] & ~x[63];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & x[15] & ~x[22] & ~x[24] & ~x[26] & ~x[27] & ~x[28] & ~x[33] & ~x[34] & ~x[35] & ~x[37] & ~x[47] & ~x[49] & ~x[50] & ~x[52] & ~x[53] & ~x[55] & ~x[58] & ~x[59] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[251] 	= partial_clause_prev[251] & ~x[0] & x[42];
			partial_clause[252] 	= partial_clause_prev[252] & ~x[2] & ~x[4] & ~x[5] & ~x[27] & ~x[30] & ~x[33] & ~x[35] & ~x[52];
			partial_clause[253] 	= partial_clause_prev[253] & 1'b1;
			partial_clause[254] 	= partial_clause_prev[254] & 1'b1;
			partial_clause[255] 	= partial_clause_prev[255] & ~x[31];
			partial_clause[256] 	= partial_clause_prev[256] & x[20];
			partial_clause[257] 	= partial_clause_prev[257] & ~x[3] & ~x[31];
			partial_clause[258] 	= partial_clause_prev[258] & ~x[23] & ~x[29] & ~x[58];
			partial_clause[259] 	= partial_clause_prev[259] & 1'b1;
			partial_clause[260] 	= partial_clause_prev[260] & ~x[9] & ~x[26] & ~x[35] & x[43] & ~x[61] & ~x[63];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[3] & ~x[4] & x[13] & ~x[24] & ~x[29] & ~x[31] & x[41] & ~x[52] & ~x[56];
			partial_clause[262] 	= partial_clause_prev[262] & ~x[60];
			partial_clause[263] 	= partial_clause_prev[263] & x[15] & ~x[26] & ~x[29] & ~x[33];
			partial_clause[264] 	= partial_clause_prev[264] & ~x[20] & ~x[25];
			partial_clause[265] 	= partial_clause_prev[265] & ~x[10] & ~x[12];
			partial_clause[266] 	= partial_clause_prev[266] & ~x[2] & ~x[6] & ~x[25] & ~x[27] & ~x[29] & ~x[35] & ~x[50] & ~x[53] & ~x[57];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[1] & ~x[25] & ~x[28] & ~x[40] & ~x[50] & ~x[52] & ~x[53] & ~x[59] & ~x[61] & ~x[62];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[2] & ~x[21] & ~x[25] & ~x[27] & ~x[30] & ~x[32] & ~x[50] & ~x[51] & ~x[54] & ~x[55] & ~x[59];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[0] & ~x[1] & ~x[2] & ~x[24] & ~x[28] & ~x[29] & ~x[30] & ~x[31] & ~x[52] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[58];
			partial_clause[270] 	= partial_clause_prev[270] & 1'b1;
			partial_clause[271] 	= partial_clause_prev[271] & ~x[13] & ~x[43] & ~x[53];
			partial_clause[272] 	= partial_clause_prev[272] & ~x[0] & ~x[1] & ~x[2] & ~x[24] & ~x[28] & ~x[59] & ~x[60];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[0] & ~x[1] & ~x[23] & ~x[25] & ~x[26] & ~x[29] & ~x[30] & ~x[32] & ~x[55] & ~x[56] & ~x[57] & ~x[59];
			partial_clause[274] 	= partial_clause_prev[274] & 1'b1;
			partial_clause[275] 	= partial_clause_prev[275] & ~x[52];
			partial_clause[276] 	= partial_clause_prev[276] & ~x[6] & ~x[9] & ~x[28] & ~x[36] & ~x[50] & ~x[56] & ~x[58];
			partial_clause[277] 	= partial_clause_prev[277] & ~x[23] & ~x[52];
			partial_clause[278] 	= partial_clause_prev[278] & 1'b1;
			partial_clause[279] 	= partial_clause_prev[279] & ~x[5] & ~x[20] & ~x[21] & ~x[29] & ~x[48] & ~x[49] & ~x[50] & ~x[55] & ~x[58] & ~x[59];
			partial_clause[280] 	= partial_clause_prev[280] & x[8] & x[36];
			partial_clause[281] 	= partial_clause_prev[281] & ~x[1] & ~x[4] & ~x[29] & ~x[55] & ~x[58];
			partial_clause[282] 	= partial_clause_prev[282] & ~x[4] & ~x[60];
			partial_clause[283] 	= partial_clause_prev[283] & x[17];
			partial_clause[284] 	= partial_clause_prev[284] & ~x[19] & ~x[22] & ~x[45];
			partial_clause[285] 	= partial_clause_prev[285] & 1'b1;
			partial_clause[286] 	= partial_clause_prev[286] & ~x[23] & ~x[38] & ~x[52];
			partial_clause[287] 	= partial_clause_prev[287] & ~x[3] & ~x[5] & ~x[21] & ~x[22] & ~x[24] & ~x[25] & ~x[26];
			partial_clause[288] 	= partial_clause_prev[288] & ~x[0] & ~x[12];
			partial_clause[289] 	= partial_clause_prev[289] & ~x[60];
			partial_clause[290] 	= partial_clause_prev[290] & ~x[1];
			partial_clause[291] 	= partial_clause_prev[291] & 1'b1;
			partial_clause[292] 	= partial_clause_prev[292] & ~x[50];
			partial_clause[293] 	= partial_clause_prev[293] & ~x[31] & ~x[33] & ~x[63];
			partial_clause[294] 	= partial_clause_prev[294] & ~x[21] & ~x[53] & ~x[60];
			partial_clause[295] 	= partial_clause_prev[295] & ~x[22] & ~x[55];
			partial_clause[296] 	= partial_clause_prev[296] & 1'b1;
			partial_clause[297] 	= partial_clause_prev[297] & ~x[24] & ~x[29] & ~x[53] & ~x[55] & ~x[63];
			partial_clause[298] 	= partial_clause_prev[298] & 1'b1;
			partial_clause[299] 	= partial_clause_prev[299] & ~x[4] & ~x[35] & ~x[50] & ~x[51] & ~x[58];
			partial_clause[300] 	= partial_clause_prev[300] & ~x[2] & ~x[5] & ~x[28];
			partial_clause[301] 	= partial_clause_prev[301] & ~x[27] & ~x[55] & ~x[62];
			partial_clause[302] 	= partial_clause_prev[302] & x[14];
			partial_clause[303] 	= partial_clause_prev[303] & ~x[38] & ~x[50];
			partial_clause[304] 	= partial_clause_prev[304] & ~x[52];
			partial_clause[305] 	= partial_clause_prev[305] & ~x[20] & ~x[31] & ~x[46] & ~x[47] & ~x[48] & ~x[50] & ~x[54] & ~x[58];
			partial_clause[306] 	= partial_clause_prev[306] & ~x[31] & ~x[61];
			partial_clause[307] 	= partial_clause_prev[307] & ~x[3] & ~x[26] & ~x[27] & ~x[28] & ~x[31] & ~x[33] & ~x[49] & ~x[59];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[0] & ~x[53] & ~x[61];
			partial_clause[309] 	= partial_clause_prev[309] & 1'b1;
			partial_clause[310] 	= partial_clause_prev[310] & ~x[50];
			partial_clause[311] 	= partial_clause_prev[311] & ~x[25] & ~x[55];
			partial_clause[312] 	= partial_clause_prev[312] & ~x[14] & ~x[51];
			partial_clause[313] 	= partial_clause_prev[313] & x[7] & ~x[52];
			partial_clause[314] 	= partial_clause_prev[314] & ~x[6] & ~x[8] & x[12] & x[39] & ~x[55] & ~x[61];
			partial_clause[315] 	= partial_clause_prev[315] & ~x[27] & ~x[30];
			partial_clause[316] 	= partial_clause_prev[316] & ~x[4] & ~x[5] & ~x[8] & ~x[10] & ~x[19] & ~x[20] & ~x[25] & ~x[27] & ~x[30] & ~x[31] & ~x[33] & ~x[37] & ~x[38] & ~x[51] & ~x[53] & ~x[54];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[24] & ~x[29] & ~x[52] & ~x[54] & ~x[58];
			partial_clause[318] 	= partial_clause_prev[318] & ~x[26] & ~x[49];
			partial_clause[319] 	= partial_clause_prev[319] & ~x[20] & ~x[51];
			partial_clause[320] 	= partial_clause_prev[320] & ~x[55] & ~x[56];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[19] & ~x[21] & ~x[23] & ~x[26] & ~x[28] & ~x[58] & ~x[59];
			partial_clause[322] 	= partial_clause_prev[322] & ~x[9] & ~x[22] & ~x[39] & ~x[41] & ~x[51];
			partial_clause[323] 	= partial_clause_prev[323] & ~x[1] & ~x[53];
			partial_clause[324] 	= partial_clause_prev[324] & ~x[41];
			partial_clause[325] 	= partial_clause_prev[325] & ~x[0] & ~x[1] & ~x[3] & ~x[24] & ~x[25] & ~x[26] & ~x[28] & ~x[56] & ~x[57];
			partial_clause[326] 	= partial_clause_prev[326] & ~x[26] & ~x[27] & ~x[28] & ~x[54] & ~x[55];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[33] & ~x[52];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[2] & ~x[57];
			partial_clause[329] 	= partial_clause_prev[329] & 1'b1;
			partial_clause[330] 	= partial_clause_prev[330] & ~x[54];
			partial_clause[331] 	= partial_clause_prev[331] & ~x[1];
			partial_clause[332] 	= partial_clause_prev[332] & ~x[2] & ~x[6] & ~x[32] & ~x[48] & ~x[50] & ~x[53] & ~x[56];
			partial_clause[333] 	= partial_clause_prev[333] & 1'b1;
			partial_clause[334] 	= partial_clause_prev[334] & ~x[29] & ~x[34];
			partial_clause[335] 	= partial_clause_prev[335] & ~x[32] & ~x[54];
			partial_clause[336] 	= partial_clause_prev[336] & ~x[41];
			partial_clause[337] 	= partial_clause_prev[337] & ~x[28];
			partial_clause[338] 	= partial_clause_prev[338] & 1'b1;
			partial_clause[339] 	= partial_clause_prev[339] & ~x[2] & ~x[8] & ~x[9] & ~x[10] & ~x[28] & ~x[31] & ~x[37] & ~x[39] & ~x[40] & ~x[52] & ~x[53];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[0] & ~x[5] & ~x[24] & ~x[50] & ~x[59] & ~x[60];
			partial_clause[341] 	= partial_clause_prev[341] & 1'b1;
			partial_clause[342] 	= partial_clause_prev[342] & ~x[0] & ~x[2] & ~x[24] & ~x[26] & ~x[58];
			partial_clause[343] 	= partial_clause_prev[343] & ~x[1] & ~x[5] & ~x[27] & ~x[61];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[24] & ~x[53];
			partial_clause[345] 	= partial_clause_prev[345] & ~x[29];
			partial_clause[346] 	= partial_clause_prev[346] & ~x[4] & ~x[5] & ~x[24] & ~x[32] & ~x[55];
			partial_clause[347] 	= partial_clause_prev[347] & ~x[0] & ~x[10] & ~x[30] & ~x[39] & ~x[40] & ~x[58];
			partial_clause[348] 	= partial_clause_prev[348] & ~x[5] & ~x[57];
			partial_clause[349] 	= partial_clause_prev[349] & ~x[29] & ~x[52] & ~x[62];
			partial_clause[350] 	= partial_clause_prev[350] & ~x[0] & ~x[1] & ~x[2] & ~x[22] & ~x[23] & ~x[25] & ~x[26] & ~x[28] & ~x[30] & ~x[31] & ~x[33] & ~x[34] & ~x[55] & ~x[57] & ~x[58];
			partial_clause[351] 	= partial_clause_prev[351] & ~x[7] & x[11] & x[39];
			partial_clause[352] 	= partial_clause_prev[352] & 1'b1;
			partial_clause[353] 	= partial_clause_prev[353] & ~x[0];
			partial_clause[354] 	= partial_clause_prev[354] & ~x[0] & ~x[1];
			partial_clause[355] 	= partial_clause_prev[355] & ~x[3] & ~x[54];
			partial_clause[356] 	= partial_clause_prev[356] & ~x[3] & ~x[10] & ~x[14] & ~x[28] & ~x[40];
			partial_clause[357] 	= partial_clause_prev[357] & 1'b1;
			partial_clause[358] 	= partial_clause_prev[358] & ~x[0] & ~x[55] & ~x[61];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[3] & ~x[4] & ~x[26] & ~x[54];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[22] & ~x[55] & ~x[61];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[33] & ~x[59] & ~x[61];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[30] & ~x[57];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[3] & ~x[4] & ~x[22] & ~x[26] & ~x[31] & ~x[50] & ~x[54] & ~x[63];
			partial_clause[364] 	= partial_clause_prev[364] & ~x[52] & ~x[55];
			partial_clause[365] 	= partial_clause_prev[365] & 1'b1;
			partial_clause[366] 	= partial_clause_prev[366] & ~x[1] & ~x[2] & ~x[4] & x[16] & ~x[29] & ~x[56] & ~x[58];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[33];
			partial_clause[368] 	= partial_clause_prev[368] & 1'b1;
			partial_clause[369] 	= partial_clause_prev[369] & x[11] & ~x[31] & ~x[53];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[2] & ~x[5] & ~x[28] & ~x[47] & ~x[49] & ~x[57];
			partial_clause[371] 	= partial_clause_prev[371] & 1'b1;
			partial_clause[372] 	= partial_clause_prev[372] & x[16] & x[17];
			partial_clause[373] 	= partial_clause_prev[373] & 1'b1;
			partial_clause[374] 	= partial_clause_prev[374] & ~x[35] & ~x[36] & ~x[55] & ~x[56];
			partial_clause[375] 	= partial_clause_prev[375] & ~x[23] & ~x[63];
			partial_clause[376] 	= partial_clause_prev[376] & ~x[1] & ~x[3] & ~x[26] & ~x[30] & ~x[31] & ~x[38] & ~x[47] & ~x[54] & ~x[60] & ~x[62];
			partial_clause[377] 	= partial_clause_prev[377] & ~x[2] & ~x[27] & ~x[28] & ~x[30];
			partial_clause[378] 	= partial_clause_prev[378] & ~x[36] & ~x[50];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[2] & ~x[33] & ~x[53] & ~x[54] & ~x[59] & ~x[60];
			partial_clause[380] 	= partial_clause_prev[380] & 1'b1;
			partial_clause[381] 	= partial_clause_prev[381] & ~x[29] & ~x[30] & ~x[32] & ~x[56] & ~x[59];
			partial_clause[382] 	= partial_clause_prev[382] & ~x[15];
			partial_clause[383] 	= partial_clause_prev[383] & 1'b1;
			partial_clause[384] 	= partial_clause_prev[384] & 1'b1;
			partial_clause[385] 	= partial_clause_prev[385] & ~x[23];
			partial_clause[386] 	= partial_clause_prev[386] & 1'b1;
			partial_clause[387] 	= partial_clause_prev[387] & ~x[2] & ~x[3] & ~x[6] & ~x[21] & ~x[22] & ~x[24] & ~x[28] & ~x[31] & ~x[33] & ~x[54] & ~x[55] & ~x[57] & ~x[58] & ~x[60] & ~x[62];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[1] & ~x[27] & ~x[31] & ~x[54] & ~x[55] & ~x[56] & ~x[58];
			partial_clause[389] 	= partial_clause_prev[389] & 1'b1;
			partial_clause[390] 	= partial_clause_prev[390] & ~x[3] & ~x[23] & ~x[24] & ~x[27] & ~x[30] & ~x[49] & ~x[50] & ~x[58];
			partial_clause[391] 	= partial_clause_prev[391] & 1'b1;
			partial_clause[392] 	= partial_clause_prev[392] & ~x[63];
			partial_clause[393] 	= partial_clause_prev[393] & 1'b1;
			partial_clause[394] 	= partial_clause_prev[394] & ~x[0];
			partial_clause[395] 	= partial_clause_prev[395] & ~x[0];
			partial_clause[396] 	= partial_clause_prev[396] & 1'b1;
			partial_clause[397] 	= partial_clause_prev[397] & 1'b1;
			partial_clause[398] 	= partial_clause_prev[398] & 1'b1;
			partial_clause[399] 	= partial_clause_prev[399] & 1'b1;
			partial_clause[400] 	= partial_clause_prev[400] & ~x[2] & ~x[4] & ~x[24] & ~x[29] & ~x[32] & ~x[34] & ~x[55] & ~x[56];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[4] & ~x[28] & ~x[32] & ~x[33] & ~x[49] & ~x[55] & ~x[56] & ~x[59];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[1] & ~x[3] & ~x[5] & ~x[7] & x[14] & ~x[23] & ~x[30] & ~x[54];
			partial_clause[403] 	= partial_clause_prev[403] & x[41];
			partial_clause[404] 	= partial_clause_prev[404] & 1'b1;
			partial_clause[405] 	= partial_clause_prev[405] & ~x[2] & ~x[3] & ~x[6] & ~x[18] & ~x[25] & ~x[51] & ~x[53];
			partial_clause[406] 	= partial_clause_prev[406] & ~x[28] & ~x[31] & ~x[57];
			partial_clause[407] 	= partial_clause_prev[407] & 1'b1;
			partial_clause[408] 	= partial_clause_prev[408] & ~x[1] & ~x[2] & ~x[21] & ~x[55];
			partial_clause[409] 	= partial_clause_prev[409] & ~x[0] & ~x[1] & ~x[5] & ~x[7] & ~x[21] & ~x[22] & ~x[25] & ~x[26] & ~x[27] & ~x[32] & ~x[51] & ~x[53] & ~x[55] & ~x[60];
			partial_clause[410] 	= partial_clause_prev[410] & x[17];
			partial_clause[411] 	= partial_clause_prev[411] & ~x[28] & x[43] & ~x[58];
			partial_clause[412] 	= partial_clause_prev[412] & ~x[1] & ~x[4] & ~x[20] & ~x[22] & ~x[25] & ~x[29] & ~x[31] & ~x[32] & ~x[52] & ~x[55];
			partial_clause[413] 	= partial_clause_prev[413] & ~x[5] & ~x[6] & ~x[18] & ~x[26] & ~x[33] & ~x[46] & ~x[47];
			partial_clause[414] 	= partial_clause_prev[414] & ~x[1] & ~x[2] & ~x[24] & ~x[25] & ~x[28] & ~x[30];
			partial_clause[415] 	= partial_clause_prev[415] & ~x[29] & ~x[58];
			partial_clause[416] 	= partial_clause_prev[416] & ~x[1] & ~x[2] & ~x[5] & ~x[23] & ~x[25] & ~x[30] & ~x[32] & ~x[49] & ~x[54] & ~x[56] & ~x[60];
			partial_clause[417] 	= partial_clause_prev[417] & ~x[0] & ~x[29] & ~x[31] & ~x[57];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[23] & ~x[30] & ~x[31] & ~x[33] & ~x[35] & ~x[49] & ~x[50] & ~x[51] & ~x[55] & ~x[57] & ~x[59];
			partial_clause[419] 	= partial_clause_prev[419] & 1'b1;
			partial_clause[420] 	= partial_clause_prev[420] & ~x[7] & x[12];
			partial_clause[421] 	= partial_clause_prev[421] & ~x[6] & ~x[22] & ~x[25] & ~x[31] & ~x[33] & ~x[55];
			partial_clause[422] 	= partial_clause_prev[422] & 1'b1;
			partial_clause[423] 	= partial_clause_prev[423] & 1'b1;
			partial_clause[424] 	= partial_clause_prev[424] & ~x[2] & ~x[18] & ~x[29] & ~x[33];
			partial_clause[425] 	= partial_clause_prev[425] & ~x[16] & ~x[25];
			partial_clause[426] 	= partial_clause_prev[426] & ~x[1] & ~x[2] & ~x[4] & ~x[5] & ~x[25] & ~x[27] & ~x[28] & ~x[30] & ~x[32] & ~x[50] & ~x[60] & ~x[63];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[0] & ~x[4] & ~x[6] & ~x[7] & ~x[27] & ~x[32] & ~x[40] & ~x[41] & ~x[50] & ~x[54];
			partial_clause[428] 	= partial_clause_prev[428] & 1'b1;
			partial_clause[429] 	= partial_clause_prev[429] & x[34];
			partial_clause[430] 	= partial_clause_prev[430] & ~x[4] & ~x[21] & ~x[23] & ~x[30] & ~x[32] & ~x[49] & ~x[51] & ~x[56] & ~x[60];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[24] & ~x[35] & ~x[36] & ~x[52];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[8] & ~x[24] & ~x[28] & ~x[29] & ~x[58];
			partial_clause[433] 	= partial_clause_prev[433] & ~x[13] & ~x[14] & ~x[27] & ~x[43] & ~x[44];
			partial_clause[434] 	= partial_clause_prev[434] & ~x[26];
			partial_clause[435] 	= partial_clause_prev[435] & ~x[0] & ~x[2] & ~x[6] & ~x[22] & ~x[34] & ~x[36] & ~x[57] & ~x[59];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[54];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[2] & ~x[26] & ~x[54] & ~x[55] & ~x[56] & ~x[57];
			partial_clause[438] 	= partial_clause_prev[438] & ~x[18] & x[43] & ~x[46] & ~x[52];
			partial_clause[439] 	= partial_clause_prev[439] & 1'b1;
			partial_clause[440] 	= partial_clause_prev[440] & ~x[33] & x[38];
			partial_clause[441] 	= partial_clause_prev[441] & 1'b1;
			partial_clause[442] 	= partial_clause_prev[442] & ~x[38];
			partial_clause[443] 	= partial_clause_prev[443] & ~x[4] & ~x[6] & ~x[29] & ~x[35] & ~x[52] & ~x[53] & ~x[55] & ~x[60] & ~x[61] & ~x[63];
			partial_clause[444] 	= partial_clause_prev[444] & ~x[40];
			partial_clause[445] 	= partial_clause_prev[445] & ~x[33];
			partial_clause[446] 	= partial_clause_prev[446] & ~x[6] & ~x[9] & ~x[29] & ~x[30] & ~x[37] & ~x[42] & ~x[54];
			partial_clause[447] 	= partial_clause_prev[447] & ~x[1] & ~x[27];
			partial_clause[448] 	= partial_clause_prev[448] & ~x[10];
			partial_clause[449] 	= partial_clause_prev[449] & ~x[25] & ~x[43] & ~x[55] & ~x[56];
			partial_clause[450] 	= partial_clause_prev[450] & ~x[26];
			partial_clause[451] 	= partial_clause_prev[451] & 1'b1;
			partial_clause[452] 	= partial_clause_prev[452] & x[14];
			partial_clause[453] 	= partial_clause_prev[453] & 1'b1;
			partial_clause[454] 	= partial_clause_prev[454] & ~x[1] & ~x[20] & ~x[47] & ~x[59];
			partial_clause[455] 	= partial_clause_prev[455] & x[15] & ~x[28] & ~x[30];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[5] & ~x[28] & ~x[49] & ~x[58] & ~x[61];
			partial_clause[457] 	= partial_clause_prev[457] & 1'b1;
			partial_clause[458] 	= partial_clause_prev[458] & ~x[10] & ~x[25] & ~x[38] & ~x[52] & ~x[54];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[25] & ~x[28];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[21] & ~x[23] & ~x[25] & ~x[26] & ~x[29] & ~x[34] & ~x[49] & ~x[55] & ~x[56];
			partial_clause[461] 	= partial_clause_prev[461] & ~x[23] & ~x[27] & ~x[29];
			partial_clause[462] 	= partial_clause_prev[462] & x[20];
			partial_clause[463] 	= partial_clause_prev[463] & x[15];
			partial_clause[464] 	= partial_clause_prev[464] & x[14] & x[15] & ~x[22] & ~x[50] & ~x[58];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[2] & ~x[3] & ~x[21] & ~x[25] & ~x[29] & ~x[30] & ~x[31] & ~x[34] & ~x[52] & ~x[53] & ~x[56];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[14] & ~x[26] & ~x[30] & ~x[42] & ~x[43] & ~x[55];
			partial_clause[467] 	= partial_clause_prev[467] & ~x[5] & ~x[7] & ~x[18] & ~x[20] & ~x[28] & ~x[45] & ~x[57];
			partial_clause[468] 	= partial_clause_prev[468] & ~x[21] & ~x[40] & ~x[54];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[5] & ~x[8] & ~x[9] & ~x[10] & ~x[28] & ~x[36] & ~x[52] & ~x[58] & ~x[63];
			partial_clause[470] 	= partial_clause_prev[470] & ~x[57];
			partial_clause[471] 	= partial_clause_prev[471] & ~x[4] & ~x[7] & ~x[23] & ~x[24] & ~x[26] & ~x[48] & ~x[51] & ~x[57] & ~x[58] & ~x[59];
			partial_clause[472] 	= partial_clause_prev[472] & 1'b1;
			partial_clause[473] 	= partial_clause_prev[473] & ~x[0] & ~x[24] & ~x[26] & ~x[28] & ~x[29] & ~x[30] & ~x[52] & ~x[53] & ~x[58];
			partial_clause[474] 	= partial_clause_prev[474] & ~x[27];
			partial_clause[475] 	= partial_clause_prev[475] & ~x[28];
			partial_clause[476] 	= partial_clause_prev[476] & 1'b1;
			partial_clause[477] 	= partial_clause_prev[477] & ~x[1] & ~x[27];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[0] & ~x[1] & ~x[25] & ~x[26] & ~x[30] & ~x[31] & ~x[32] & ~x[55] & ~x[59];
			partial_clause[479] 	= partial_clause_prev[479] & 1'b1;
			partial_clause[480] 	= partial_clause_prev[480] & ~x[0] & ~x[2] & ~x[3] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[22] & ~x[23] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[35] & ~x[49] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[59] & ~x[60];
			partial_clause[481] 	= partial_clause_prev[481] & 1'b1;
			partial_clause[482] 	= partial_clause_prev[482] & ~x[50];
			partial_clause[483] 	= partial_clause_prev[483] & 1'b1;
			partial_clause[484] 	= partial_clause_prev[484] & ~x[26] & ~x[32] & ~x[49];
			partial_clause[485] 	= partial_clause_prev[485] & 1'b1;
			partial_clause[486] 	= partial_clause_prev[486] & ~x[1] & ~x[57];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[29] & ~x[54];
			partial_clause[488] 	= partial_clause_prev[488] & 1'b1;
			partial_clause[489] 	= partial_clause_prev[489] & x[15];
			partial_clause[490] 	= partial_clause_prev[490] & ~x[46];
			partial_clause[491] 	= partial_clause_prev[491] & 1'b1;
			partial_clause[492] 	= partial_clause_prev[492] & ~x[55] & ~x[58];
			partial_clause[493] 	= partial_clause_prev[493] & x[14];
			partial_clause[494] 	= partial_clause_prev[494] & ~x[28] & ~x[60];
			partial_clause[495] 	= partial_clause_prev[495] & ~x[0] & ~x[2] & ~x[6] & ~x[7] & ~x[35] & ~x[36] & ~x[38] & ~x[56];
			partial_clause[496] 	= partial_clause_prev[496] & 1'b1;
			partial_clause[497] 	= partial_clause_prev[497] & ~x[0] & ~x[10] & ~x[11] & ~x[27] & ~x[63];
			partial_clause[498] 	= partial_clause_prev[498] & 1'b1;
			partial_clause[499] 	= partial_clause_prev[499] & 1'b1;
		end
	end
endmodule


module HCB_8 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[18] & ~x[20] & ~x[22] & ~x[45] & ~x[48] & ~x[50];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[12] & ~x[13] & ~x[25] & ~x[38] & ~x[53];
			partial_clause[2] 	= partial_clause_prev[2] & ~x[2] & ~x[4] & ~x[20];
			partial_clause[3] 	= partial_clause_prev[3] & ~x[15];
			partial_clause[4] 	= partial_clause_prev[4] & ~x[45];
			partial_clause[5] 	= partial_clause_prev[5] & ~x[15] & ~x[22] & ~x[48];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[16];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[20] & ~x[52];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[17] & ~x[21] & ~x[22] & ~x[50];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[2] & ~x[5] & ~x[16] & ~x[17] & ~x[31] & ~x[47] & ~x[50] & ~x[51];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[15] & ~x[16] & ~x[24] & ~x[42] & ~x[47] & ~x[52];
			partial_clause[11] 	= partial_clause_prev[11] & x[8] & x[9] & ~x[13] & x[35] & ~x[43] & ~x[48] & ~x[49];
			partial_clause[12] 	= partial_clause_prev[12] & ~x[44] & ~x[45] & ~x[46] & ~x[48];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[10] & ~x[14] & ~x[15] & ~x[20] & ~x[22] & ~x[38] & ~x[39] & ~x[41] & ~x[43] & ~x[49] & ~x[51];
			partial_clause[14] 	= partial_clause_prev[14] & 1'b1;
			partial_clause[15] 	= partial_clause_prev[15] & 1'b1;
			partial_clause[16] 	= partial_clause_prev[16] & ~x[16] & ~x[17] & ~x[18] & ~x[22] & ~x[23];
			partial_clause[17] 	= partial_clause_prev[17] & 1'b1;
			partial_clause[18] 	= partial_clause_prev[18] & ~x[21];
			partial_clause[19] 	= partial_clause_prev[19] & ~x[4] & ~x[6] & ~x[7] & ~x[45] & ~x[49] & ~x[50] & ~x[53];
			partial_clause[20] 	= partial_clause_prev[20] & 1'b1;
			partial_clause[21] 	= partial_clause_prev[21] & 1'b1;
			partial_clause[22] 	= partial_clause_prev[22] & ~x[40] & ~x[42] & ~x[44] & ~x[48];
			partial_clause[23] 	= partial_clause_prev[23] & ~x[18] & ~x[19] & ~x[47] & ~x[48] & ~x[49];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[17] & ~x[18] & ~x[20] & ~x[48] & ~x[49] & ~x[50] & ~x[52] & ~x[54];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[12] & ~x[14] & ~x[23] & ~x[24] & ~x[25] & ~x[38] & ~x[43] & ~x[46] & ~x[47] & ~x[50] & ~x[52];
			partial_clause[26] 	= partial_clause_prev[26] & ~x[4];
			partial_clause[27] 	= partial_clause_prev[27] & ~x[18] & ~x[21] & ~x[22];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[17] & ~x[38];
			partial_clause[29] 	= partial_clause_prev[29] & ~x[25] & ~x[45];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[5] & ~x[19];
			partial_clause[31] 	= partial_clause_prev[31] & 1'b1;
			partial_clause[32] 	= partial_clause_prev[32] & ~x[12] & ~x[51];
			partial_clause[33] 	= partial_clause_prev[33] & 1'b1;
			partial_clause[34] 	= partial_clause_prev[34] & ~x[14] & ~x[18] & ~x[20] & ~x[21] & ~x[22] & ~x[24] & ~x[46] & ~x[50];
			partial_clause[35] 	= partial_clause_prev[35] & ~x[16] & ~x[17] & ~x[19] & ~x[44] & ~x[45];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[19];
			partial_clause[37] 	= partial_clause_prev[37] & ~x[22] & ~x[48] & ~x[58];
			partial_clause[38] 	= partial_clause_prev[38] & ~x[15] & ~x[18] & ~x[20] & ~x[21];
			partial_clause[39] 	= partial_clause_prev[39] & ~x[38];
			partial_clause[40] 	= partial_clause_prev[40] & ~x[18] & ~x[19] & ~x[31];
			partial_clause[41] 	= partial_clause_prev[41] & x[2];
			partial_clause[42] 	= partial_clause_prev[42] & 1'b1;
			partial_clause[43] 	= partial_clause_prev[43] & ~x[21] & ~x[47];
			partial_clause[44] 	= partial_clause_prev[44] & 1'b1;
			partial_clause[45] 	= partial_clause_prev[45] & 1'b1;
			partial_clause[46] 	= partial_clause_prev[46] & ~x[19] & ~x[21] & ~x[44] & ~x[45] & ~x[54];
			partial_clause[47] 	= partial_clause_prev[47] & ~x[27] & ~x[28];
			partial_clause[48] 	= partial_clause_prev[48] & 1'b1;
			partial_clause[49] 	= partial_clause_prev[49] & 1'b1;
			partial_clause[50] 	= partial_clause_prev[50] & ~x[24] & x[30] & x[58];
			partial_clause[51] 	= partial_clause_prev[51] & 1'b1;
			partial_clause[52] 	= partial_clause_prev[52] & 1'b1;
			partial_clause[53] 	= partial_clause_prev[53] & 1'b1;
			partial_clause[54] 	= partial_clause_prev[54] & ~x[58];
			partial_clause[55] 	= partial_clause_prev[55] & 1'b1;
			partial_clause[56] 	= partial_clause_prev[56] & 1'b1;
			partial_clause[57] 	= partial_clause_prev[57] & ~x[18];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[17] & ~x[21] & ~x[39] & ~x[40] & ~x[42];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[14] & ~x[24] & ~x[25] & ~x[42] & ~x[46] & ~x[47] & ~x[51] & ~x[59] & ~x[60];
			partial_clause[60] 	= partial_clause_prev[60] & ~x[2] & ~x[3] & ~x[6] & ~x[32];
			partial_clause[61] 	= partial_clause_prev[61] & 1'b1;
			partial_clause[62] 	= partial_clause_prev[62] & ~x[3] & ~x[13] & ~x[14] & ~x[15] & ~x[30] & ~x[45];
			partial_clause[63] 	= partial_clause_prev[63] & ~x[18] & ~x[47];
			partial_clause[64] 	= partial_clause_prev[64] & ~x[47];
			partial_clause[65] 	= partial_clause_prev[65] & x[33];
			partial_clause[66] 	= partial_clause_prev[66] & 1'b1;
			partial_clause[67] 	= partial_clause_prev[67] & 1'b1;
			partial_clause[68] 	= partial_clause_prev[68] & ~x[48];
			partial_clause[69] 	= partial_clause_prev[69] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[21] & ~x[32] & ~x[43] & ~x[46] & ~x[49] & ~x[51];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[16];
			partial_clause[71] 	= partial_clause_prev[71] & ~x[2] & ~x[4];
			partial_clause[72] 	= partial_clause_prev[72] & 1'b1;
			partial_clause[73] 	= partial_clause_prev[73] & ~x[25];
			partial_clause[74] 	= partial_clause_prev[74] & ~x[17] & ~x[20] & ~x[21];
			partial_clause[75] 	= partial_clause_prev[75] & 1'b1;
			partial_clause[76] 	= partial_clause_prev[76] & ~x[13] & ~x[16] & ~x[18] & ~x[20] & ~x[21] & ~x[25] & ~x[41] & ~x[45] & ~x[50] & ~x[52];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[46];
			partial_clause[78] 	= partial_clause_prev[78] & ~x[53];
			partial_clause[79] 	= partial_clause_prev[79] & ~x[0] & ~x[15] & ~x[37] & ~x[41] & ~x[44];
			partial_clause[80] 	= partial_clause_prev[80] & 1'b1;
			partial_clause[81] 	= partial_clause_prev[81] & x[3] & ~x[18] & x[30];
			partial_clause[82] 	= partial_clause_prev[82] & ~x[49];
			partial_clause[83] 	= partial_clause_prev[83] & x[4] & x[31];
			partial_clause[84] 	= partial_clause_prev[84] & ~x[1];
			partial_clause[85] 	= partial_clause_prev[85] & ~x[13] & ~x[17] & ~x[58];
			partial_clause[86] 	= partial_clause_prev[86] & x[4] & ~x[27] & ~x[28] & x[32] & ~x[42];
			partial_clause[87] 	= partial_clause_prev[87] & 1'b1;
			partial_clause[88] 	= partial_clause_prev[88] & ~x[5] & ~x[6] & ~x[17] & ~x[46];
			partial_clause[89] 	= partial_clause_prev[89] & ~x[23];
			partial_clause[90] 	= partial_clause_prev[90] & ~x[57];
			partial_clause[91] 	= partial_clause_prev[91] & 1'b1;
			partial_clause[92] 	= partial_clause_prev[92] & ~x[19] & ~x[41] & ~x[42] & ~x[49];
			partial_clause[93] 	= partial_clause_prev[93] & ~x[18] & ~x[19] & ~x[47] & ~x[48] & ~x[53] & ~x[54];
			partial_clause[94] 	= partial_clause_prev[94] & 1'b1;
			partial_clause[95] 	= partial_clause_prev[95] & ~x[17] & ~x[19] & ~x[23] & ~x[24] & ~x[27] & ~x[45];
			partial_clause[96] 	= partial_clause_prev[96] & ~x[31];
			partial_clause[97] 	= partial_clause_prev[97] & ~x[14] & ~x[23] & ~x[41] & ~x[42] & ~x[47] & ~x[53];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[19] & ~x[45] & ~x[49] & ~x[50] & ~x[51] & ~x[52];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[15] & ~x[18] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[26] & ~x[42] & ~x[43] & ~x[46] & ~x[48] & ~x[49] & ~x[52] & ~x[53] & ~x[54];
			partial_clause[100] 	= partial_clause_prev[100] & ~x[19];
			partial_clause[101] 	= partial_clause_prev[101] & ~x[33];
			partial_clause[102] 	= partial_clause_prev[102] & ~x[11] & ~x[12] & ~x[40];
			partial_clause[103] 	= partial_clause_prev[103] & ~x[14] & ~x[17] & ~x[18] & ~x[21] & ~x[22] & ~x[41] & ~x[49];
			partial_clause[104] 	= partial_clause_prev[104] & 1'b1;
			partial_clause[105] 	= partial_clause_prev[105] & ~x[2] & ~x[13] & ~x[16] & ~x[17] & ~x[19] & ~x[20] & ~x[24] & ~x[26] & ~x[31] & ~x[38] & ~x[40] & ~x[42] & ~x[53] & ~x[54] & ~x[58];
			partial_clause[106] 	= partial_clause_prev[106] & ~x[24];
			partial_clause[107] 	= partial_clause_prev[107] & ~x[14] & ~x[16] & ~x[17] & ~x[21] & ~x[26] & ~x[38] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[47] & ~x[53] & ~x[54] & ~x[55] & ~x[56];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[25] & ~x[29] & ~x[46] & ~x[47] & ~x[54];
			partial_clause[109] 	= partial_clause_prev[109] & 1'b1;
			partial_clause[110] 	= partial_clause_prev[110] & x[6] & ~x[44] & x[62];
			partial_clause[111] 	= partial_clause_prev[111] & 1'b1;
			partial_clause[112] 	= partial_clause_prev[112] & ~x[6] & ~x[49];
			partial_clause[113] 	= partial_clause_prev[113] & 1'b1;
			partial_clause[114] 	= partial_clause_prev[114] & x[25];
			partial_clause[115] 	= partial_clause_prev[115] & ~x[15] & ~x[16] & ~x[17] & ~x[19] & ~x[22] & ~x[34] & ~x[46] & ~x[48] & ~x[51] & ~x[53] & ~x[55];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[12] & ~x[18] & ~x[20] & ~x[24];
			partial_clause[117] 	= partial_clause_prev[117] & 1'b1;
			partial_clause[118] 	= partial_clause_prev[118] & ~x[1] & ~x[19];
			partial_clause[119] 	= partial_clause_prev[119] & ~x[16] & ~x[18] & ~x[20] & ~x[21] & ~x[22] & ~x[26] & ~x[31] & ~x[32] & ~x[43] & ~x[48] & ~x[49] & ~x[54] & ~x[56] & ~x[59] & ~x[60];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[17] & ~x[18] & ~x[19] & ~x[21] & ~x[35] & ~x[45] & ~x[46] & ~x[47] & ~x[49] & ~x[51] & ~x[52];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[18] & ~x[22] & x[38];
			partial_clause[122] 	= partial_clause_prev[122] & ~x[11];
			partial_clause[123] 	= partial_clause_prev[123] & ~x[15] & ~x[16] & ~x[17] & ~x[21] & ~x[23] & ~x[51];
			partial_clause[124] 	= partial_clause_prev[124] & x[59];
			partial_clause[125] 	= partial_clause_prev[125] & ~x[22] & ~x[23] & ~x[24];
			partial_clause[126] 	= partial_clause_prev[126] & ~x[12] & ~x[41] & ~x[45] & ~x[53] & ~x[55];
			partial_clause[127] 	= partial_clause_prev[127] & ~x[21] & ~x[24] & ~x[25] & ~x[26] & ~x[43] & ~x[44] & ~x[47] & ~x[50] & ~x[51];
			partial_clause[128] 	= partial_clause_prev[128] & ~x[22];
			partial_clause[129] 	= partial_clause_prev[129] & ~x[19] & ~x[24] & ~x[25];
			partial_clause[130] 	= partial_clause_prev[130] & 1'b1;
			partial_clause[131] 	= partial_clause_prev[131] & ~x[15] & ~x[27];
			partial_clause[132] 	= partial_clause_prev[132] & ~x[55] & ~x[56];
			partial_clause[133] 	= partial_clause_prev[133] & ~x[12] & ~x[24] & ~x[29] & ~x[38] & ~x[46];
			partial_clause[134] 	= partial_clause_prev[134] & ~x[18] & ~x[19] & ~x[21] & ~x[23] & ~x[42] & ~x[48] & ~x[49];
			partial_clause[135] 	= partial_clause_prev[135] & ~x[42];
			partial_clause[136] 	= partial_clause_prev[136] & ~x[14] & ~x[16] & ~x[43] & ~x[44] & ~x[45];
			partial_clause[137] 	= partial_clause_prev[137] & ~x[29];
			partial_clause[138] 	= partial_clause_prev[138] & ~x[0] & ~x[1] & ~x[3];
			partial_clause[139] 	= partial_clause_prev[139] & ~x[15] & ~x[22] & ~x[23] & ~x[47] & ~x[48] & ~x[50];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[18] & ~x[21] & ~x[42] & ~x[47] & ~x[48] & ~x[49];
			partial_clause[141] 	= partial_clause_prev[141] & ~x[3] & ~x[4] & ~x[16];
			partial_clause[142] 	= partial_clause_prev[142] & ~x[19] & ~x[21] & ~x[25] & ~x[28] & ~x[43] & ~x[46] & ~x[47] & ~x[48] & ~x[52] & ~x[53] & ~x[54];
			partial_clause[143] 	= partial_clause_prev[143] & ~x[20];
			partial_clause[144] 	= partial_clause_prev[144] & ~x[14] & ~x[16] & ~x[19] & ~x[46];
			partial_clause[145] 	= partial_clause_prev[145] & 1'b1;
			partial_clause[146] 	= partial_clause_prev[146] & ~x[12] & ~x[13] & ~x[18] & ~x[20] & ~x[39] & ~x[40];
			partial_clause[147] 	= partial_clause_prev[147] & ~x[14] & ~x[24] & ~x[50] & ~x[52];
			partial_clause[148] 	= partial_clause_prev[148] & x[7] & ~x[16] & ~x[20] & ~x[25] & ~x[41] & ~x[43] & ~x[54] & ~x[55] & ~x[56] & ~x[59];
			partial_clause[149] 	= partial_clause_prev[149] & ~x[24];
			partial_clause[150] 	= partial_clause_prev[150] & ~x[14] & ~x[21] & ~x[22];
			partial_clause[151] 	= partial_clause_prev[151] & ~x[8];
			partial_clause[152] 	= partial_clause_prev[152] & ~x[14] & ~x[57];
			partial_clause[153] 	= partial_clause_prev[153] & ~x[3] & ~x[5] & ~x[7] & ~x[18] & ~x[24] & ~x[29] & ~x[46] & ~x[47] & ~x[51] & ~x[52];
			partial_clause[154] 	= partial_clause_prev[154] & 1'b1;
			partial_clause[155] 	= partial_clause_prev[155] & 1'b1;
			partial_clause[156] 	= partial_clause_prev[156] & x[31];
			partial_clause[157] 	= partial_clause_prev[157] & 1'b1;
			partial_clause[158] 	= partial_clause_prev[158] & ~x[11] & ~x[16] & ~x[22] & ~x[24] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[50];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[16] & ~x[19] & ~x[23] & ~x[26] & ~x[52];
			partial_clause[160] 	= partial_clause_prev[160] & ~x[11] & ~x[15] & ~x[47] & ~x[50];
			partial_clause[161] 	= partial_clause_prev[161] & ~x[14] & ~x[21] & ~x[26] & ~x[28] & ~x[29] & ~x[42] & ~x[43] & ~x[46] & ~x[48];
			partial_clause[162] 	= partial_clause_prev[162] & ~x[19] & ~x[46] & ~x[49] & ~x[50];
			partial_clause[163] 	= partial_clause_prev[163] & 1'b1;
			partial_clause[164] 	= partial_clause_prev[164] & ~x[39];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[29] & ~x[42] & ~x[43] & ~x[47] & ~x[55] & ~x[57];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[24] & ~x[51] & x[57];
			partial_clause[167] 	= partial_clause_prev[167] & 1'b1;
			partial_clause[168] 	= partial_clause_prev[168] & ~x[22];
			partial_clause[169] 	= partial_clause_prev[169] & ~x[18] & ~x[23] & ~x[53];
			partial_clause[170] 	= partial_clause_prev[170] & 1'b1;
			partial_clause[171] 	= partial_clause_prev[171] & ~x[18] & ~x[19] & ~x[49] & ~x[53];
			partial_clause[172] 	= partial_clause_prev[172] & 1'b1;
			partial_clause[173] 	= partial_clause_prev[173] & ~x[17] & ~x[44];
			partial_clause[174] 	= partial_clause_prev[174] & ~x[16] & ~x[37] & ~x[38] & ~x[40] & ~x[45] & ~x[53];
			partial_clause[175] 	= partial_clause_prev[175] & 1'b1;
			partial_clause[176] 	= partial_clause_prev[176] & ~x[50];
			partial_clause[177] 	= partial_clause_prev[177] & ~x[39] & ~x[53];
			partial_clause[178] 	= partial_clause_prev[178] & ~x[53];
			partial_clause[179] 	= partial_clause_prev[179] & 1'b1;
			partial_clause[180] 	= partial_clause_prev[180] & ~x[1] & ~x[16] & ~x[25] & ~x[31] & ~x[33];
			partial_clause[181] 	= partial_clause_prev[181] & x[1] & x[28] & x[56];
			partial_clause[182] 	= partial_clause_prev[182] & ~x[15];
			partial_clause[183] 	= partial_clause_prev[183] & ~x[2] & ~x[3] & ~x[19] & ~x[45] & ~x[49] & ~x[51];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[11] & ~x[12] & ~x[13] & ~x[28] & ~x[41] & ~x[45] & ~x[51];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[16] & ~x[19] & ~x[50] & x[61];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[11] & ~x[22] & ~x[24] & ~x[44] & ~x[48] & ~x[51] & ~x[53];
			partial_clause[187] 	= partial_clause_prev[187] & ~x[15] & ~x[21] & ~x[24] & ~x[44] & ~x[50] & ~x[60] & ~x[61];
			partial_clause[188] 	= partial_clause_prev[188] & 1'b1;
			partial_clause[189] 	= partial_clause_prev[189] & ~x[3];
			partial_clause[190] 	= partial_clause_prev[190] & ~x[11] & ~x[12] & ~x[14] & ~x[17] & ~x[25] & ~x[55] & ~x[57];
			partial_clause[191] 	= partial_clause_prev[191] & ~x[22];
			partial_clause[192] 	= partial_clause_prev[192] & ~x[5] & ~x[7] & ~x[48] & ~x[51];
			partial_clause[193] 	= partial_clause_prev[193] & ~x[17] & ~x[54];
			partial_clause[194] 	= partial_clause_prev[194] & 1'b1;
			partial_clause[195] 	= partial_clause_prev[195] & ~x[10] & ~x[14] & ~x[21] & ~x[22] & ~x[44] & ~x[54];
			partial_clause[196] 	= partial_clause_prev[196] & ~x[21];
			partial_clause[197] 	= partial_clause_prev[197] & ~x[15] & ~x[21] & ~x[48];
			partial_clause[198] 	= partial_clause_prev[198] & ~x[24];
			partial_clause[199] 	= partial_clause_prev[199] & x[27];
			partial_clause[200] 	= partial_clause_prev[200] & ~x[2] & ~x[3] & ~x[6] & ~x[9] & ~x[23] & ~x[34] & ~x[50];
			partial_clause[201] 	= partial_clause_prev[201] & ~x[22] & ~x[41] & ~x[43];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[17] & ~x[19] & ~x[44] & ~x[47] & ~x[52];
			partial_clause[203] 	= partial_clause_prev[203] & ~x[12] & ~x[16] & ~x[42];
			partial_clause[204] 	= partial_clause_prev[204] & ~x[1] & ~x[14] & ~x[18] & ~x[22] & ~x[25] & ~x[27] & ~x[41] & ~x[43] & ~x[46] & ~x[53];
			partial_clause[205] 	= partial_clause_prev[205] & 1'b1;
			partial_clause[206] 	= partial_clause_prev[206] & ~x[16] & ~x[17] & ~x[20] & ~x[44];
			partial_clause[207] 	= partial_clause_prev[207] & ~x[23] & ~x[40];
			partial_clause[208] 	= partial_clause_prev[208] & ~x[16] & ~x[17] & ~x[30] & ~x[42] & ~x[43];
			partial_clause[209] 	= partial_clause_prev[209] & x[33] & x[60];
			partial_clause[210] 	= partial_clause_prev[210] & ~x[19] & ~x[22] & ~x[41] & ~x[42];
			partial_clause[211] 	= partial_clause_prev[211] & ~x[11] & ~x[15];
			partial_clause[212] 	= partial_clause_prev[212] & ~x[18] & ~x[42];
			partial_clause[213] 	= partial_clause_prev[213] & 1'b1;
			partial_clause[214] 	= partial_clause_prev[214] & ~x[19];
			partial_clause[215] 	= partial_clause_prev[215] & x[1] & ~x[23];
			partial_clause[216] 	= partial_clause_prev[216] & ~x[15];
			partial_clause[217] 	= partial_clause_prev[217] & ~x[18] & ~x[23] & ~x[51];
			partial_clause[218] 	= partial_clause_prev[218] & 1'b1;
			partial_clause[219] 	= partial_clause_prev[219] & 1'b1;
			partial_clause[220] 	= partial_clause_prev[220] & ~x[12] & ~x[16] & ~x[18] & ~x[40] & ~x[45] & ~x[46] & ~x[48];
			partial_clause[221] 	= partial_clause_prev[221] & ~x[2] & ~x[29] & ~x[46] & ~x[55];
			partial_clause[222] 	= partial_clause_prev[222] & 1'b1;
			partial_clause[223] 	= partial_clause_prev[223] & ~x[36] & ~x[54];
			partial_clause[224] 	= partial_clause_prev[224] & ~x[14] & ~x[15] & ~x[16] & ~x[33] & ~x[48] & ~x[60];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[44] & ~x[49];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[14] & ~x[22] & ~x[44] & ~x[49] & ~x[53];
			partial_clause[227] 	= partial_clause_prev[227] & x[5] & x[31];
			partial_clause[228] 	= partial_clause_prev[228] & ~x[11] & ~x[13] & ~x[17] & ~x[19] & ~x[22] & ~x[44] & ~x[47];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[16] & ~x[17] & ~x[24] & ~x[48] & ~x[51] & ~x[52];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[14] & ~x[15] & ~x[18] & ~x[19] & ~x[22] & ~x[23] & ~x[41] & ~x[43] & ~x[44] & ~x[47] & ~x[49];
			partial_clause[231] 	= partial_clause_prev[231] & ~x[16] & ~x[17] & ~x[46] & ~x[47];
			partial_clause[232] 	= partial_clause_prev[232] & 1'b1;
			partial_clause[233] 	= partial_clause_prev[233] & ~x[17];
			partial_clause[234] 	= partial_clause_prev[234] & ~x[22];
			partial_clause[235] 	= partial_clause_prev[235] & 1'b1;
			partial_clause[236] 	= partial_clause_prev[236] & x[8] & ~x[39] & ~x[41];
			partial_clause[237] 	= partial_clause_prev[237] & ~x[15];
			partial_clause[238] 	= partial_clause_prev[238] & ~x[9] & ~x[39] & ~x[48];
			partial_clause[239] 	= partial_clause_prev[239] & x[32];
			partial_clause[240] 	= partial_clause_prev[240] & ~x[18] & ~x[22] & ~x[45] & ~x[50];
			partial_clause[241] 	= partial_clause_prev[241] & ~x[16] & ~x[23] & ~x[54];
			partial_clause[242] 	= partial_clause_prev[242] & ~x[14] & ~x[19] & ~x[21] & ~x[22] & ~x[42] & ~x[47] & ~x[52];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[17] & ~x[18] & ~x[19] & ~x[23] & ~x[47] & ~x[50] & ~x[51];
			partial_clause[244] 	= partial_clause_prev[244] & ~x[30] & ~x[31] & ~x[47] & ~x[58] & ~x[59];
			partial_clause[245] 	= partial_clause_prev[245] & 1'b1;
			partial_clause[246] 	= partial_clause_prev[246] & ~x[18] & ~x[48];
			partial_clause[247] 	= partial_clause_prev[247] & ~x[13] & ~x[14] & ~x[20] & ~x[21] & ~x[24] & ~x[26] & ~x[41] & ~x[44] & ~x[47] & ~x[50] & ~x[51];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[15] & ~x[20] & ~x[43] & ~x[54];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[4] & ~x[16];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[0] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[20] & ~x[22] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & ~x[39] & ~x[41] & ~x[44] & ~x[47] & ~x[48] & ~x[50] & ~x[52];
			partial_clause[251] 	= partial_clause_prev[251] & ~x[37];
			partial_clause[252] 	= partial_clause_prev[252] & ~x[18] & ~x[23] & ~x[24] & ~x[44] & ~x[47] & ~x[51] & ~x[53] & ~x[54];
			partial_clause[253] 	= partial_clause_prev[253] & ~x[52];
			partial_clause[254] 	= partial_clause_prev[254] & ~x[16];
			partial_clause[255] 	= partial_clause_prev[255] & ~x[23] & ~x[24] & x[35];
			partial_clause[256] 	= partial_clause_prev[256] & 1'b1;
			partial_clause[257] 	= partial_clause_prev[257] & ~x[31] & ~x[44] & ~x[47];
			partial_clause[258] 	= partial_clause_prev[258] & ~x[16] & ~x[24] & ~x[43] & ~x[45] & ~x[51] & ~x[52] & ~x[58];
			partial_clause[259] 	= partial_clause_prev[259] & 1'b1;
			partial_clause[260] 	= partial_clause_prev[260] & ~x[17] & ~x[48] & ~x[53];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[20] & ~x[41] & ~x[46] & ~x[47] & ~x[52];
			partial_clause[262] 	= partial_clause_prev[262] & 1'b1;
			partial_clause[263] 	= partial_clause_prev[263] & ~x[16];
			partial_clause[264] 	= partial_clause_prev[264] & ~x[17] & ~x[40] & ~x[41];
			partial_clause[265] 	= partial_clause_prev[265] & 1'b1;
			partial_clause[266] 	= partial_clause_prev[266] & ~x[14] & ~x[17] & ~x[20] & ~x[21] & ~x[44] & ~x[49] & ~x[54];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[3] & ~x[4] & ~x[18] & ~x[19] & ~x[20] & ~x[26] & ~x[27] & ~x[43] & ~x[49] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[54] & ~x[55];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[13] & ~x[14] & ~x[20] & ~x[22] & ~x[30] & ~x[42] & ~x[44] & ~x[49] & ~x[50];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[18] & ~x[22] & ~x[43] & ~x[44] & ~x[45] & ~x[47] & ~x[48] & ~x[51] & ~x[52];
			partial_clause[270] 	= partial_clause_prev[270] & 1'b1;
			partial_clause[271] 	= partial_clause_prev[271] & 1'b1;
			partial_clause[272] 	= partial_clause_prev[272] & ~x[48];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[16] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[45] & ~x[48] & ~x[50] & ~x[52] & ~x[53] & ~x[54];
			partial_clause[274] 	= partial_clause_prev[274] & ~x[50];
			partial_clause[275] 	= partial_clause_prev[275] & ~x[49] & ~x[58];
			partial_clause[276] 	= partial_clause_prev[276] & ~x[23] & ~x[47] & ~x[48] & ~x[51] & ~x[53] & ~x[55];
			partial_clause[277] 	= partial_clause_prev[277] & ~x[17] & ~x[24] & ~x[54];
			partial_clause[278] 	= partial_clause_prev[278] & ~x[6];
			partial_clause[279] 	= partial_clause_prev[279] & ~x[11] & ~x[15] & ~x[16] & ~x[17] & ~x[23] & ~x[40] & ~x[43] & ~x[44] & ~x[46] & ~x[48] & ~x[51] & ~x[52];
			partial_clause[280] 	= partial_clause_prev[280] & 1'b1;
			partial_clause[281] 	= partial_clause_prev[281] & 1'b1;
			partial_clause[282] 	= partial_clause_prev[282] & x[57];
			partial_clause[283] 	= partial_clause_prev[283] & ~x[21];
			partial_clause[284] 	= partial_clause_prev[284] & 1'b1;
			partial_clause[285] 	= partial_clause_prev[285] & 1'b1;
			partial_clause[286] 	= partial_clause_prev[286] & ~x[37] & ~x[50];
			partial_clause[287] 	= partial_clause_prev[287] & ~x[6] & ~x[15] & ~x[18] & ~x[44] & ~x[46] & ~x[51];
			partial_clause[288] 	= partial_clause_prev[288] & 1'b1;
			partial_clause[289] 	= partial_clause_prev[289] & ~x[20] & ~x[47];
			partial_clause[290] 	= partial_clause_prev[290] & 1'b1;
			partial_clause[291] 	= partial_clause_prev[291] & ~x[42];
			partial_clause[292] 	= partial_clause_prev[292] & ~x[17] & ~x[21] & ~x[54];
			partial_clause[293] 	= partial_clause_prev[293] & ~x[16] & ~x[19] & ~x[52] & ~x[54];
			partial_clause[294] 	= partial_clause_prev[294] & ~x[52];
			partial_clause[295] 	= partial_clause_prev[295] & 1'b1;
			partial_clause[296] 	= partial_clause_prev[296] & 1'b1;
			partial_clause[297] 	= partial_clause_prev[297] & ~x[28] & ~x[29] & ~x[41] & ~x[44] & ~x[52] & ~x[54];
			partial_clause[298] 	= partial_clause_prev[298] & 1'b1;
			partial_clause[299] 	= partial_clause_prev[299] & ~x[43] & ~x[52];
			partial_clause[300] 	= partial_clause_prev[300] & ~x[17] & ~x[23];
			partial_clause[301] 	= partial_clause_prev[301] & ~x[12] & ~x[15] & ~x[28] & ~x[40] & ~x[58];
			partial_clause[302] 	= partial_clause_prev[302] & ~x[25] & ~x[28];
			partial_clause[303] 	= partial_clause_prev[303] & ~x[1] & ~x[13] & ~x[24] & ~x[46];
			partial_clause[304] 	= partial_clause_prev[304] & ~x[17];
			partial_clause[305] 	= partial_clause_prev[305] & ~x[7] & ~x[34] & ~x[62];
			partial_clause[306] 	= partial_clause_prev[306] & ~x[50] & ~x[52];
			partial_clause[307] 	= partial_clause_prev[307] & ~x[15] & ~x[17] & ~x[23] & ~x[26] & ~x[27] & ~x[40] & ~x[49] & ~x[55];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[16] & ~x[22];
			partial_clause[309] 	= partial_clause_prev[309] & ~x[23] & ~x[51];
			partial_clause[310] 	= partial_clause_prev[310] & 1'b1;
			partial_clause[311] 	= partial_clause_prev[311] & ~x[28] & ~x[46] & ~x[56] & ~x[63];
			partial_clause[312] 	= partial_clause_prev[312] & ~x[16] & ~x[42];
			partial_clause[313] 	= partial_clause_prev[313] & ~x[17];
			partial_clause[314] 	= partial_clause_prev[314] & x[2] & ~x[51];
			partial_clause[315] 	= partial_clause_prev[315] & ~x[18] & ~x[28] & ~x[29] & ~x[41] & ~x[43];
			partial_clause[316] 	= partial_clause_prev[316] & ~x[0] & ~x[2] & ~x[14] & ~x[21] & ~x[27] & ~x[44] & ~x[47] & ~x[50];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[17] & ~x[46] & ~x[57];
			partial_clause[318] 	= partial_clause_prev[318] & ~x[18];
			partial_clause[319] 	= partial_clause_prev[319] & ~x[11];
			partial_clause[320] 	= partial_clause_prev[320] & ~x[17] & ~x[46] & ~x[48];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[13] & ~x[17] & ~x[20] & ~x[25] & ~x[40] & ~x[41] & ~x[43] & ~x[45] & ~x[48] & ~x[51];
			partial_clause[322] 	= partial_clause_prev[322] & ~x[16] & ~x[21] & ~x[42] & ~x[45] & ~x[48];
			partial_clause[323] 	= partial_clause_prev[323] & ~x[13] & ~x[22] & ~x[25] & ~x[57];
			partial_clause[324] 	= partial_clause_prev[324] & ~x[3] & ~x[4] & ~x[5];
			partial_clause[325] 	= partial_clause_prev[325] & ~x[13] & ~x[18] & ~x[21] & ~x[23] & ~x[42] & ~x[43] & ~x[49];
			partial_clause[326] 	= partial_clause_prev[326] & ~x[20] & ~x[47];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[27] & ~x[43] & ~x[45] & ~x[46] & x[62] & x[63];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[22] & ~x[23];
			partial_clause[329] 	= partial_clause_prev[329] & 1'b1;
			partial_clause[330] 	= partial_clause_prev[330] & x[3] & ~x[45];
			partial_clause[331] 	= partial_clause_prev[331] & ~x[12];
			partial_clause[332] 	= partial_clause_prev[332] & ~x[26] & ~x[48] & ~x[51];
			partial_clause[333] 	= partial_clause_prev[333] & 1'b1;
			partial_clause[334] 	= partial_clause_prev[334] & ~x[17];
			partial_clause[335] 	= partial_clause_prev[335] & ~x[16];
			partial_clause[336] 	= partial_clause_prev[336] & 1'b1;
			partial_clause[337] 	= partial_clause_prev[337] & 1'b1;
			partial_clause[338] 	= partial_clause_prev[338] & x[61];
			partial_clause[339] 	= partial_clause_prev[339] & ~x[4] & ~x[16] & ~x[21] & ~x[23] & ~x[51];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[19] & ~x[26] & ~x[43] & ~x[45] & ~x[47] & ~x[49] & ~x[52] & ~x[58] & ~x[59];
			partial_clause[341] 	= partial_clause_prev[341] & 1'b1;
			partial_clause[342] 	= partial_clause_prev[342] & ~x[17] & ~x[19] & ~x[50];
			partial_clause[343] 	= partial_clause_prev[343] & ~x[17] & ~x[20] & ~x[21] & ~x[22] & ~x[45] & ~x[51];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[42] & ~x[47];
			partial_clause[345] 	= partial_clause_prev[345] & 1'b1;
			partial_clause[346] 	= partial_clause_prev[346] & ~x[20];
			partial_clause[347] 	= partial_clause_prev[347] & ~x[4] & ~x[5] & ~x[16] & ~x[51];
			partial_clause[348] 	= partial_clause_prev[348] & ~x[18] & ~x[36];
			partial_clause[349] 	= partial_clause_prev[349] & ~x[43] & ~x[48] & ~x[52];
			partial_clause[350] 	= partial_clause_prev[350] & ~x[18] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[47] & ~x[48] & ~x[49] & ~x[51] & ~x[54];
			partial_clause[351] 	= partial_clause_prev[351] & ~x[24];
			partial_clause[352] 	= partial_clause_prev[352] & 1'b1;
			partial_clause[353] 	= partial_clause_prev[353] & ~x[59];
			partial_clause[354] 	= partial_clause_prev[354] & ~x[19];
			partial_clause[355] 	= partial_clause_prev[355] & ~x[48];
			partial_clause[356] 	= partial_clause_prev[356] & ~x[45] & ~x[48];
			partial_clause[357] 	= partial_clause_prev[357] & x[12] & x[40];
			partial_clause[358] 	= partial_clause_prev[358] & ~x[11] & ~x[19] & ~x[21] & ~x[41] & ~x[52] & ~x[56];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[47] & ~x[50];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[4] & ~x[16] & ~x[21] & ~x[22] & ~x[23] & ~x[27] & ~x[29] & ~x[31] & ~x[42] & ~x[43] & ~x[48] & ~x[50] & ~x[53] & ~x[56] & ~x[58] & ~x[59];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[18] & ~x[23] & ~x[44] & ~x[48] & ~x[49];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[21] & ~x[49] & ~x[51] & ~x[63];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[24] & ~x[26] & ~x[39] & ~x[40] & ~x[43] & ~x[48] & ~x[51] & ~x[52] & ~x[53];
			partial_clause[364] 	= partial_clause_prev[364] & ~x[14] & ~x[21] & ~x[49];
			partial_clause[365] 	= partial_clause_prev[365] & 1'b1;
			partial_clause[366] 	= partial_clause_prev[366] & ~x[15] & ~x[17] & ~x[20] & ~x[22] & ~x[24] & ~x[41] & ~x[42] & ~x[46] & ~x[49] & ~x[50] & ~x[52] & ~x[55];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[43];
			partial_clause[368] 	= partial_clause_prev[368] & 1'b1;
			partial_clause[369] 	= partial_clause_prev[369] & ~x[16] & ~x[23] & ~x[27] & ~x[30] & ~x[31] & ~x[56];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[11] & ~x[12] & ~x[16] & ~x[21] & ~x[37] & ~x[40] & ~x[41] & ~x[50] & ~x[54];
			partial_clause[371] 	= partial_clause_prev[371] & 1'b1;
			partial_clause[372] 	= partial_clause_prev[372] & ~x[26] & ~x[27] & ~x[50] & ~x[55];
			partial_clause[373] 	= partial_clause_prev[373] & 1'b1;
			partial_clause[374] 	= partial_clause_prev[374] & ~x[2] & ~x[3] & ~x[18] & ~x[20] & ~x[24] & ~x[33] & ~x[34];
			partial_clause[375] 	= partial_clause_prev[375] & ~x[45];
			partial_clause[376] 	= partial_clause_prev[376] & ~x[2] & ~x[11] & ~x[12] & ~x[16] & ~x[30] & ~x[44] & ~x[47] & ~x[49] & ~x[57];
			partial_clause[377] 	= partial_clause_prev[377] & ~x[47];
			partial_clause[378] 	= partial_clause_prev[378] & ~x[3] & ~x[43];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[21];
			partial_clause[380] 	= partial_clause_prev[380] & 1'b1;
			partial_clause[381] 	= partial_clause_prev[381] & ~x[22];
			partial_clause[382] 	= partial_clause_prev[382] & 1'b1;
			partial_clause[383] 	= partial_clause_prev[383] & 1'b1;
			partial_clause[384] 	= partial_clause_prev[384] & 1'b1;
			partial_clause[385] 	= partial_clause_prev[385] & 1'b1;
			partial_clause[386] 	= partial_clause_prev[386] & 1'b1;
			partial_clause[387] 	= partial_clause_prev[387] & ~x[17] & ~x[18] & ~x[23] & ~x[47] & ~x[48] & ~x[50];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[17] & ~x[18] & ~x[19] & ~x[22] & ~x[24] & ~x[40] & ~x[47] & ~x[48] & ~x[50] & ~x[51];
			partial_clause[389] 	= partial_clause_prev[389] & 1'b1;
			partial_clause[390] 	= partial_clause_prev[390] & ~x[13] & ~x[18] & ~x[19] & ~x[43] & ~x[44];
			partial_clause[391] 	= partial_clause_prev[391] & 1'b1;
			partial_clause[392] 	= partial_clause_prev[392] & ~x[35] & ~x[63];
			partial_clause[393] 	= partial_clause_prev[393] & 1'b1;
			partial_clause[394] 	= partial_clause_prev[394] & 1'b1;
			partial_clause[395] 	= partial_clause_prev[395] & x[38];
			partial_clause[396] 	= partial_clause_prev[396] & x[13];
			partial_clause[397] 	= partial_clause_prev[397] & 1'b1;
			partial_clause[398] 	= partial_clause_prev[398] & ~x[4];
			partial_clause[399] 	= partial_clause_prev[399] & 1'b1;
			partial_clause[400] 	= partial_clause_prev[400] & ~x[42] & ~x[47] & ~x[48] & ~x[51] & ~x[52];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[13] & ~x[45] & ~x[46] & ~x[52];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[14] & ~x[15] & ~x[18] & ~x[19] & ~x[21] & ~x[24] & ~x[42] & ~x[49];
			partial_clause[403] 	= partial_clause_prev[403] & ~x[24] & ~x[28] & ~x[53] & ~x[57] & x[60];
			partial_clause[404] 	= partial_clause_prev[404] & x[31];
			partial_clause[405] 	= partial_clause_prev[405] & ~x[41] & ~x[43] & ~x[47];
			partial_clause[406] 	= partial_clause_prev[406] & x[9] & ~x[24];
			partial_clause[407] 	= partial_clause_prev[407] & ~x[16];
			partial_clause[408] 	= partial_clause_prev[408] & ~x[14] & ~x[18];
			partial_clause[409] 	= partial_clause_prev[409] & ~x[15] & ~x[19] & ~x[20] & ~x[22] & ~x[23] & ~x[24] & ~x[42] & ~x[45] & ~x[51] & ~x[52] & ~x[53] & ~x[55];
			partial_clause[410] 	= partial_clause_prev[410] & ~x[50] & ~x[58];
			partial_clause[411] 	= partial_clause_prev[411] & 1'b1;
			partial_clause[412] 	= partial_clause_prev[412] & ~x[16] & ~x[23] & ~x[25] & ~x[42] & ~x[46] & ~x[50];
			partial_clause[413] 	= partial_clause_prev[413] & ~x[19];
			partial_clause[414] 	= partial_clause_prev[414] & ~x[17] & ~x[19] & ~x[21] & ~x[23] & ~x[43] & ~x[45] & ~x[51];
			partial_clause[415] 	= partial_clause_prev[415] & ~x[21] & ~x[24] & ~x[48] & ~x[52];
			partial_clause[416] 	= partial_clause_prev[416] & ~x[15] & ~x[23] & ~x[41] & ~x[51];
			partial_clause[417] 	= partial_clause_prev[417] & ~x[17] & ~x[32] & ~x[48];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[0] & ~x[12] & ~x[16] & ~x[17] & ~x[20] & ~x[21] & ~x[22] & ~x[24] & ~x[29] & ~x[41] & ~x[46] & ~x[52];
			partial_clause[419] 	= partial_clause_prev[419] & 1'b1;
			partial_clause[420] 	= partial_clause_prev[420] & x[61];
			partial_clause[421] 	= partial_clause_prev[421] & ~x[23] & ~x[52] & ~x[53];
			partial_clause[422] 	= partial_clause_prev[422] & ~x[14] & ~x[43] & ~x[50];
			partial_clause[423] 	= partial_clause_prev[423] & ~x[20] & x[41] & ~x[49];
			partial_clause[424] 	= partial_clause_prev[424] & 1'b1;
			partial_clause[425] 	= partial_clause_prev[425] & ~x[19];
			partial_clause[426] 	= partial_clause_prev[426] & ~x[14] & ~x[16] & ~x[19] & ~x[46] & ~x[48] & ~x[51];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[2] & ~x[5] & ~x[29] & ~x[44] & ~x[46] & ~x[47];
			partial_clause[428] 	= partial_clause_prev[428] & 1'b1;
			partial_clause[429] 	= partial_clause_prev[429] & 1'b1;
			partial_clause[430] 	= partial_clause_prev[430] & ~x[15] & ~x[16] & ~x[24] & ~x[39] & ~x[50] & ~x[52];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[2] & ~x[19];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[17] & ~x[20] & ~x[23] & ~x[45];
			partial_clause[433] 	= partial_clause_prev[433] & ~x[19] & ~x[20];
			partial_clause[434] 	= partial_clause_prev[434] & ~x[23] & ~x[32] & ~x[54] & ~x[57];
			partial_clause[435] 	= partial_clause_prev[435] & ~x[13] & ~x[15] & ~x[19] & ~x[20] & ~x[22] & ~x[23] & ~x[41] & ~x[42] & ~x[45] & ~x[48] & ~x[51];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[18] & ~x[21];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[18] & ~x[24] & ~x[41] & ~x[42] & ~x[44] & ~x[51];
			partial_clause[438] 	= partial_clause_prev[438] & 1'b1;
			partial_clause[439] 	= partial_clause_prev[439] & ~x[20];
			partial_clause[440] 	= partial_clause_prev[440] & x[30] & ~x[50];
			partial_clause[441] 	= partial_clause_prev[441] & ~x[17] & ~x[22] & ~x[46];
			partial_clause[442] 	= partial_clause_prev[442] & ~x[27];
			partial_clause[443] 	= partial_clause_prev[443] & ~x[17] & ~x[19] & ~x[24] & ~x[25] & ~x[26] & ~x[28] & ~x[46] & ~x[49];
			partial_clause[444] 	= partial_clause_prev[444] & 1'b1;
			partial_clause[445] 	= partial_clause_prev[445] & ~x[38];
			partial_clause[446] 	= partial_clause_prev[446] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[33] & ~x[43] & ~x[45] & ~x[47] & ~x[48];
			partial_clause[447] 	= partial_clause_prev[447] & ~x[20] & ~x[21] & ~x[23] & ~x[48];
			partial_clause[448] 	= partial_clause_prev[448] & 1'b1;
			partial_clause[449] 	= partial_clause_prev[449] & ~x[19] & ~x[50] & ~x[51] & ~x[53];
			partial_clause[450] 	= partial_clause_prev[450] & ~x[1] & ~x[11] & ~x[14] & ~x[24] & ~x[27] & ~x[31] & ~x[43] & ~x[47];
			partial_clause[451] 	= partial_clause_prev[451] & x[61];
			partial_clause[452] 	= partial_clause_prev[452] & ~x[48];
			partial_clause[453] 	= partial_clause_prev[453] & ~x[33] & ~x[57];
			partial_clause[454] 	= partial_clause_prev[454] & ~x[39] & ~x[48];
			partial_clause[455] 	= partial_clause_prev[455] & ~x[18] & ~x[44] & ~x[57];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[16] & ~x[17] & ~x[21] & ~x[22] & ~x[24] & ~x[43] & ~x[48] & ~x[51];
			partial_clause[457] 	= partial_clause_prev[457] & 1'b1;
			partial_clause[458] 	= partial_clause_prev[458] & ~x[18] & ~x[19] & ~x[21] & ~x[45] & ~x[50];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[18];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[18] & ~x[40] & ~x[43] & ~x[50];
			partial_clause[461] 	= partial_clause_prev[461] & ~x[16] & ~x[23] & ~x[43] & ~x[49] & ~x[58] & ~x[60];
			partial_clause[462] 	= partial_clause_prev[462] & ~x[20];
			partial_clause[463] 	= partial_clause_prev[463] & 1'b1;
			partial_clause[464] 	= partial_clause_prev[464] & ~x[25] & ~x[27] & ~x[52] & ~x[53];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[19] & ~x[20] & ~x[24] & ~x[49] & ~x[53];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[18] & ~x[49] & ~x[50];
			partial_clause[467] 	= partial_clause_prev[467] & ~x[24];
			partial_clause[468] 	= partial_clause_prev[468] & ~x[42];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[15] & ~x[24] & ~x[45] & ~x[49] & ~x[55];
			partial_clause[470] 	= partial_clause_prev[470] & 1'b1;
			partial_clause[471] 	= partial_clause_prev[471] & ~x[18] & ~x[40];
			partial_clause[472] 	= partial_clause_prev[472] & ~x[16] & ~x[24] & ~x[42];
			partial_clause[473] 	= partial_clause_prev[473] & ~x[6] & ~x[16] & ~x[44] & ~x[45] & ~x[50];
			partial_clause[474] 	= partial_clause_prev[474] & ~x[35] & ~x[62];
			partial_clause[475] 	= partial_clause_prev[475] & ~x[16] & ~x[18] & ~x[23] & ~x[41] & ~x[53];
			partial_clause[476] 	= partial_clause_prev[476] & ~x[48];
			partial_clause[477] 	= partial_clause_prev[477] & ~x[18] & ~x[46];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[17] & ~x[19] & ~x[22] & ~x[24] & ~x[45] & ~x[51] & ~x[52];
			partial_clause[479] 	= partial_clause_prev[479] & x[58];
			partial_clause[480] 	= partial_clause_prev[480] & ~x[14] & ~x[15] & ~x[16] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[23] & ~x[42] & ~x[43] & ~x[45] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[52];
			partial_clause[481] 	= partial_clause_prev[481] & ~x[49];
			partial_clause[482] 	= partial_clause_prev[482] & ~x[15] & ~x[21] & ~x[41] & ~x[51];
			partial_clause[483] 	= partial_clause_prev[483] & x[8] & ~x[14];
			partial_clause[484] 	= partial_clause_prev[484] & 1'b1;
			partial_clause[485] 	= partial_clause_prev[485] & 1'b1;
			partial_clause[486] 	= partial_clause_prev[486] & ~x[48];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[23] & ~x[52];
			partial_clause[488] 	= partial_clause_prev[488] & ~x[1];
			partial_clause[489] 	= partial_clause_prev[489] & ~x[20];
			partial_clause[490] 	= partial_clause_prev[490] & 1'b1;
			partial_clause[491] 	= partial_clause_prev[491] & x[6] & ~x[22];
			partial_clause[492] 	= partial_clause_prev[492] & 1'b1;
			partial_clause[493] 	= partial_clause_prev[493] & ~x[15] & ~x[46];
			partial_clause[494] 	= partial_clause_prev[494] & ~x[18] & ~x[47];
			partial_clause[495] 	= partial_clause_prev[495] & ~x[3] & ~x[5] & ~x[6] & ~x[21] & ~x[24] & ~x[30] & ~x[32] & ~x[34] & ~x[51];
			partial_clause[496] 	= partial_clause_prev[496] & ~x[32];
			partial_clause[497] 	= partial_clause_prev[497] & ~x[46];
			partial_clause[498] 	= partial_clause_prev[498] & 1'b1;
			partial_clause[499] 	= partial_clause_prev[499] & ~x[48];
		end
	end
endmodule


module HCB_9 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[10] & ~x[11] & ~x[13] & ~x[14] & ~x[33] & ~x[36] & ~x[38] & ~x[39] & ~x[40] & ~x[42] & ~x[62] & ~x[63];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[35] & ~x[37] & ~x[41] & ~x[62];
			partial_clause[2] 	= partial_clause_prev[2] & 1'b1;
			partial_clause[3] 	= partial_clause_prev[3] & ~x[3] & ~x[40];
			partial_clause[4] 	= partial_clause_prev[4] & ~x[6] & ~x[10] & ~x[41];
			partial_clause[5] 	= partial_clause_prev[5] & ~x[7] & ~x[9] & ~x[14] & ~x[42];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[14] & x[52];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[7] & ~x[9] & ~x[18] & ~x[36] & ~x[37] & ~x[40] & ~x[46];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[4] & ~x[6] & ~x[9] & ~x[11] & ~x[14] & ~x[36] & ~x[38] & ~x[42] & ~x[58] & ~x[61];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[34] & ~x[37] & ~x[43] & ~x[44];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[4] & ~x[5] & ~x[10] & ~x[15] & ~x[40] & ~x[43] & ~x[44] & ~x[60] & ~x[62];
			partial_clause[11] 	= partial_clause_prev[11] & ~x[6] & ~x[9] & ~x[37] & ~x[61];
			partial_clause[12] 	= partial_clause_prev[12] & ~x[38] & ~x[40] & ~x[45];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[8] & ~x[31] & ~x[33] & ~x[38] & ~x[40] & ~x[43] & ~x[58] & ~x[59] & ~x[60] & ~x[61];
			partial_clause[14] 	= partial_clause_prev[14] & 1'b1;
			partial_clause[15] 	= partial_clause_prev[15] & 1'b1;
			partial_clause[16] 	= partial_clause_prev[16] & ~x[6] & ~x[14] & ~x[32] & ~x[39] & ~x[43] & ~x[60];
			partial_clause[17] 	= partial_clause_prev[17] & 1'b1;
			partial_clause[18] 	= partial_clause_prev[18] & ~x[34];
			partial_clause[19] 	= partial_clause_prev[19] & ~x[13] & ~x[40] & ~x[62] & ~x[63];
			partial_clause[20] 	= partial_clause_prev[20] & ~x[23] & ~x[24] & ~x[37] & ~x[46] & ~x[50];
			partial_clause[21] 	= partial_clause_prev[21] & ~x[13] & ~x[34] & ~x[60];
			partial_clause[22] 	= partial_clause_prev[22] & 1'b1;
			partial_clause[23] 	= partial_clause_prev[23] & ~x[9] & ~x[10] & ~x[11] & ~x[13] & ~x[14] & ~x[39] & ~x[41] & ~x[42];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[8] & ~x[10] & ~x[11] & ~x[12] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[35] & ~x[37] & ~x[38] & ~x[39] & ~x[40] & ~x[41] & ~x[44] & ~x[61] & ~x[63];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[4] & ~x[7] & ~x[8] & ~x[14] & ~x[32] & ~x[40] & ~x[41] & ~x[45];
			partial_clause[26] 	= partial_clause_prev[26] & 1'b1;
			partial_clause[27] 	= partial_clause_prev[27] & ~x[39] & ~x[42];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[1] & ~x[2] & ~x[9] & ~x[63];
			partial_clause[29] 	= partial_clause_prev[29] & ~x[9] & ~x[12] & ~x[13] & ~x[41] & ~x[44] & ~x[45];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[36];
			partial_clause[31] 	= partial_clause_prev[31] & ~x[40] & ~x[42] & ~x[43];
			partial_clause[32] 	= partial_clause_prev[32] & ~x[10] & ~x[38];
			partial_clause[33] 	= partial_clause_prev[33] & 1'b1;
			partial_clause[34] 	= partial_clause_prev[34] & ~x[8] & ~x[39];
			partial_clause[35] 	= partial_clause_prev[35] & ~x[8] & ~x[35] & ~x[36];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[14] & ~x[37] & ~x[40] & ~x[41] & ~x[63];
			partial_clause[37] 	= partial_clause_prev[37] & ~x[22] & ~x[44];
			partial_clause[38] 	= partial_clause_prev[38] & ~x[14] & x[24] & x[25] & ~x[41] & ~x[43];
			partial_clause[39] 	= partial_clause_prev[39] & ~x[2] & ~x[29] & ~x[59];
			partial_clause[40] 	= partial_clause_prev[40] & ~x[62];
			partial_clause[41] 	= partial_clause_prev[41] & ~x[48];
			partial_clause[42] 	= partial_clause_prev[42] & 1'b1;
			partial_clause[43] 	= partial_clause_prev[43] & ~x[12] & x[29] & ~x[44];
			partial_clause[44] 	= partial_clause_prev[44] & 1'b1;
			partial_clause[45] 	= partial_clause_prev[45] & ~x[9];
			partial_clause[46] 	= partial_clause_prev[46] & ~x[6] & ~x[11] & ~x[13] & ~x[14] & ~x[16] & ~x[31] & ~x[37] & ~x[40] & ~x[58] & ~x[60] & ~x[62];
			partial_clause[47] 	= partial_clause_prev[47] & ~x[3] & ~x[7] & ~x[17] & ~x[31] & ~x[44];
			partial_clause[48] 	= partial_clause_prev[48] & 1'b1;
			partial_clause[49] 	= partial_clause_prev[49] & ~x[39];
			partial_clause[50] 	= partial_clause_prev[50] & ~x[15] & ~x[43];
			partial_clause[51] 	= partial_clause_prev[51] & 1'b1;
			partial_clause[52] 	= partial_clause_prev[52] & ~x[16];
			partial_clause[53] 	= partial_clause_prev[53] & 1'b1;
			partial_clause[54] 	= partial_clause_prev[54] & ~x[6] & ~x[21] & ~x[46];
			partial_clause[55] 	= partial_clause_prev[55] & ~x[35] & ~x[61];
			partial_clause[56] 	= partial_clause_prev[56] & 1'b1;
			partial_clause[57] 	= partial_clause_prev[57] & ~x[39] & ~x[43] & ~x[46];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[4] & ~x[8] & ~x[31] & ~x[58] & ~x[61];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[10] & ~x[13] & ~x[14] & ~x[16] & ~x[17] & ~x[18] & ~x[33] & ~x[37] & ~x[41] & ~x[43] & ~x[44] & ~x[46];
			partial_clause[60] 	= partial_clause_prev[60] & ~x[63];
			partial_clause[61] 	= partial_clause_prev[61] & 1'b1;
			partial_clause[62] 	= partial_clause_prev[62] & ~x[7] & ~x[10] & ~x[11] & ~x[22] & ~x[39] & ~x[40] & ~x[46] & ~x[47] & ~x[61] & ~x[62];
			partial_clause[63] 	= partial_clause_prev[63] & 1'b1;
			partial_clause[64] 	= partial_clause_prev[64] & ~x[8];
			partial_clause[65] 	= partial_clause_prev[65] & 1'b1;
			partial_clause[66] 	= partial_clause_prev[66] & 1'b1;
			partial_clause[67] 	= partial_clause_prev[67] & ~x[62];
			partial_clause[68] 	= partial_clause_prev[68] & ~x[6] & ~x[13] & ~x[32];
			partial_clause[69] 	= partial_clause_prev[69] & ~x[42];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[42];
			partial_clause[71] 	= partial_clause_prev[71] & 1'b1;
			partial_clause[72] 	= partial_clause_prev[72] & ~x[5] & ~x[30] & ~x[41] & ~x[43] & ~x[58] & ~x[60];
			partial_clause[73] 	= partial_clause_prev[73] & 1'b1;
			partial_clause[74] 	= partial_clause_prev[74] & ~x[13];
			partial_clause[75] 	= partial_clause_prev[75] & ~x[61] & ~x[63];
			partial_clause[76] 	= partial_clause_prev[76] & ~x[5] & ~x[7] & ~x[17] & ~x[34] & ~x[37] & ~x[43] & ~x[63];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[16];
			partial_clause[78] 	= partial_clause_prev[78] & 1'b1;
			partial_clause[79] 	= partial_clause_prev[79] & ~x[2] & ~x[12] & ~x[14] & ~x[29] & ~x[58];
			partial_clause[80] 	= partial_clause_prev[80] & ~x[48];
			partial_clause[81] 	= partial_clause_prev[81] & ~x[40];
			partial_clause[82] 	= partial_clause_prev[82] & ~x[60];
			partial_clause[83] 	= partial_clause_prev[83] & 1'b1;
			partial_clause[84] 	= partial_clause_prev[84] & ~x[17] & ~x[35];
			partial_clause[85] 	= partial_clause_prev[85] & ~x[4] & ~x[16] & ~x[18] & ~x[32] & ~x[34] & ~x[41] & ~x[62];
			partial_clause[86] 	= partial_clause_prev[86] & ~x[11] & ~x[13] & ~x[15] & ~x[16] & ~x[18] & ~x[45] & ~x[47] & ~x[61] & ~x[63];
			partial_clause[87] 	= partial_clause_prev[87] & 1'b1;
			partial_clause[88] 	= partial_clause_prev[88] & ~x[8] & ~x[43];
			partial_clause[89] 	= partial_clause_prev[89] & ~x[8];
			partial_clause[90] 	= partial_clause_prev[90] & ~x[20];
			partial_clause[91] 	= partial_clause_prev[91] & ~x[60] & ~x[63];
			partial_clause[92] 	= partial_clause_prev[92] & ~x[3] & ~x[13];
			partial_clause[93] 	= partial_clause_prev[93] & ~x[9] & ~x[10] & ~x[12] & ~x[15] & ~x[18] & ~x[34] & ~x[39] & ~x[40] & ~x[45] & ~x[46] & ~x[61];
			partial_clause[94] 	= partial_clause_prev[94] & 1'b1;
			partial_clause[95] 	= partial_clause_prev[95] & ~x[6] & ~x[17] & ~x[34] & ~x[36] & ~x[41] & ~x[48] & ~x[62];
			partial_clause[96] 	= partial_clause_prev[96] & 1'b1;
			partial_clause[97] 	= partial_clause_prev[97] & ~x[5] & ~x[10] & ~x[15] & ~x[16] & ~x[33] & ~x[37] & ~x[38] & ~x[40] & ~x[61];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[10] & ~x[17] & x[23] & ~x[36] & ~x[37] & ~x[43] & x[53];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[6] & ~x[7] & ~x[9] & ~x[11] & ~x[12] & ~x[13] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[35] & ~x[39] & ~x[42] & ~x[43] & ~x[44] & ~x[46] & ~x[63];
			partial_clause[100] 	= partial_clause_prev[100] & ~x[15];
			partial_clause[101] 	= partial_clause_prev[101] & 1'b1;
			partial_clause[102] 	= partial_clause_prev[102] & 1'b1;
			partial_clause[103] 	= partial_clause_prev[103] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[11] & ~x[14] & ~x[16] & ~x[32] & ~x[33] & ~x[38] & ~x[40] & ~x[42] & ~x[43] & ~x[44] & ~x[59] & ~x[60];
			partial_clause[104] 	= partial_clause_prev[104] & ~x[14] & ~x[15] & ~x[32] & ~x[58];
			partial_clause[105] 	= partial_clause_prev[105] & ~x[8] & ~x[15] & ~x[19] & ~x[21] & ~x[30] & ~x[31] & ~x[35] & ~x[37] & ~x[39] & ~x[42] & ~x[46] & ~x[49] & ~x[60] & ~x[63];
			partial_clause[106] 	= partial_clause_prev[106] & ~x[14] & ~x[36] & ~x[40];
			partial_clause[107] 	= partial_clause_prev[107] & ~x[2] & ~x[6] & ~x[7] & ~x[10] & ~x[17] & ~x[19] & ~x[44] & ~x[45] & ~x[46] & ~x[47] & ~x[58] & ~x[59] & ~x[63];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[12] & ~x[15] & ~x[21] & ~x[36] & ~x[41] & ~x[48];
			partial_clause[109] 	= partial_clause_prev[109] & 1'b1;
			partial_clause[110] 	= partial_clause_prev[110] & ~x[51];
			partial_clause[111] 	= partial_clause_prev[111] & 1'b1;
			partial_clause[112] 	= partial_clause_prev[112] & ~x[15] & ~x[36];
			partial_clause[113] 	= partial_clause_prev[113] & ~x[4] & ~x[13] & ~x[14] & ~x[30] & ~x[37];
			partial_clause[114] 	= partial_clause_prev[114] & 1'b1;
			partial_clause[115] 	= partial_clause_prev[115] & ~x[8] & ~x[9] & ~x[11] & ~x[13] & ~x[14] & ~x[16] & ~x[36] & ~x[41] & ~x[45] & ~x[46];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[45] & ~x[62];
			partial_clause[117] 	= partial_clause_prev[117] & ~x[8];
			partial_clause[118] 	= partial_clause_prev[118] & ~x[8] & ~x[10] & ~x[20] & ~x[37];
			partial_clause[119] 	= partial_clause_prev[119] & ~x[4] & ~x[7] & ~x[10] & ~x[22] & ~x[40] & ~x[42];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[9] & ~x[11] & ~x[15] & ~x[16] & ~x[38] & ~x[40] & ~x[41] & ~x[42] & ~x[44] & x[52];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[11] & ~x[38] & ~x[39];
			partial_clause[122] 	= partial_clause_prev[122] & ~x[2] & ~x[3];
			partial_clause[123] 	= partial_clause_prev[123] & ~x[7] & ~x[11] & ~x[34] & ~x[36] & ~x[39] & ~x[40] & ~x[41] & ~x[43] & ~x[62];
			partial_clause[124] 	= partial_clause_prev[124] & 1'b1;
			partial_clause[125] 	= partial_clause_prev[125] & 1'b1;
			partial_clause[126] 	= partial_clause_prev[126] & ~x[34];
			partial_clause[127] 	= partial_clause_prev[127] & ~x[6] & ~x[8] & ~x[10] & ~x[12] & ~x[16] & ~x[17] & ~x[37] & ~x[38] & ~x[42] & ~x[43] & ~x[45] & ~x[46] & ~x[63];
			partial_clause[128] 	= partial_clause_prev[128] & ~x[45] & ~x[46];
			partial_clause[129] 	= partial_clause_prev[129] & ~x[6] & ~x[7] & ~x[12] & ~x[31] & ~x[36] & ~x[40] & ~x[61];
			partial_clause[130] 	= partial_clause_prev[130] & ~x[8] & ~x[18] & ~x[39] & ~x[40] & ~x[42] & ~x[43];
			partial_clause[131] 	= partial_clause_prev[131] & ~x[23] & ~x[44] & ~x[49] & ~x[50] & ~x[58];
			partial_clause[132] 	= partial_clause_prev[132] & ~x[14] & ~x[16] & ~x[34] & ~x[44] & ~x[47];
			partial_clause[133] 	= partial_clause_prev[133] & ~x[37] & ~x[56];
			partial_clause[134] 	= partial_clause_prev[134] & ~x[9] & ~x[11] & ~x[13] & ~x[35] & ~x[37] & ~x[38] & ~x[41] & ~x[61] & ~x[63];
			partial_clause[135] 	= partial_clause_prev[135] & x[19] & ~x[44] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[136] 	= partial_clause_prev[136] & ~x[6] & ~x[13] & ~x[32] & ~x[38] & ~x[62];
			partial_clause[137] 	= partial_clause_prev[137] & ~x[19];
			partial_clause[138] 	= partial_clause_prev[138] & x[21];
			partial_clause[139] 	= partial_clause_prev[139] & ~x[8] & ~x[10] & ~x[14] & ~x[15] & ~x[18] & ~x[37] & ~x[40] & ~x[42] & ~x[46];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[12] & ~x[15] & ~x[34] & ~x[36] & ~x[38] & ~x[40] & ~x[41] & ~x[63];
			partial_clause[141] 	= partial_clause_prev[141] & ~x[17] & ~x[23] & ~x[36] & ~x[44] & ~x[51] & ~x[62];
			partial_clause[142] 	= partial_clause_prev[142] & ~x[10] & ~x[18] & ~x[32] & ~x[33] & ~x[37] & ~x[42] & ~x[60];
			partial_clause[143] 	= partial_clause_prev[143] & 1'b1;
			partial_clause[144] 	= partial_clause_prev[144] & ~x[10] & ~x[34] & ~x[41] & ~x[42] & ~x[44] & ~x[45] & ~x[62] & ~x[63];
			partial_clause[145] 	= partial_clause_prev[145] & ~x[8];
			partial_clause[146] 	= partial_clause_prev[146] & ~x[11] & ~x[15] & ~x[16] & ~x[33] & ~x[37] & ~x[39] & ~x[60] & ~x[62];
			partial_clause[147] 	= partial_clause_prev[147] & ~x[6] & ~x[15] & ~x[16] & ~x[17] & ~x[36] & ~x[39] & ~x[41] & ~x[45] & ~x[62];
			partial_clause[148] 	= partial_clause_prev[148] & ~x[3] & ~x[4] & ~x[7] & ~x[18] & ~x[48] & ~x[62];
			partial_clause[149] 	= partial_clause_prev[149] & ~x[63];
			partial_clause[150] 	= partial_clause_prev[150] & ~x[6] & ~x[11] & ~x[35] & ~x[36] & ~x[38] & ~x[40] & ~x[42];
			partial_clause[151] 	= partial_clause_prev[151] & ~x[55];
			partial_clause[152] 	= partial_clause_prev[152] & ~x[37];
			partial_clause[153] 	= partial_clause_prev[153] & ~x[11] & ~x[14] & ~x[40];
			partial_clause[154] 	= partial_clause_prev[154] & 1'b1;
			partial_clause[155] 	= partial_clause_prev[155] & 1'b1;
			partial_clause[156] 	= partial_clause_prev[156] & 1'b1;
			partial_clause[157] 	= partial_clause_prev[157] & 1'b1;
			partial_clause[158] 	= partial_clause_prev[158] & ~x[5] & ~x[8] & ~x[10] & ~x[11] & ~x[12] & ~x[32] & ~x[35] & ~x[37] & ~x[41] & ~x[42] & ~x[59];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[9];
			partial_clause[160] 	= partial_clause_prev[160] & ~x[11] & ~x[44];
			partial_clause[161] 	= partial_clause_prev[161] & ~x[9] & ~x[10] & ~x[11] & ~x[16] & ~x[34] & ~x[36] & ~x[39] & ~x[63];
			partial_clause[162] 	= partial_clause_prev[162] & ~x[11] & ~x[16] & ~x[33] & ~x[60] & ~x[61];
			partial_clause[163] 	= partial_clause_prev[163] & 1'b1;
			partial_clause[164] 	= partial_clause_prev[164] & ~x[30] & ~x[58];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[2] & ~x[7] & ~x[12] & ~x[17] & ~x[31] & ~x[32] & ~x[39] & ~x[43] & ~x[44] & ~x[47] & ~x[62];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[9] & ~x[12] & ~x[13] & ~x[41];
			partial_clause[167] 	= partial_clause_prev[167] & 1'b1;
			partial_clause[168] 	= partial_clause_prev[168] & ~x[17] & ~x[25];
			partial_clause[169] 	= partial_clause_prev[169] & 1'b1;
			partial_clause[170] 	= partial_clause_prev[170] & ~x[49];
			partial_clause[171] 	= partial_clause_prev[171] & ~x[6] & ~x[12] & ~x[37] & ~x[42];
			partial_clause[172] 	= partial_clause_prev[172] & 1'b1;
			partial_clause[173] 	= partial_clause_prev[173] & ~x[32] & ~x[39] & ~x[62];
			partial_clause[174] 	= partial_clause_prev[174] & ~x[6] & ~x[39] & ~x[45];
			partial_clause[175] 	= partial_clause_prev[175] & 1'b1;
			partial_clause[176] 	= partial_clause_prev[176] & 1'b1;
			partial_clause[177] 	= partial_clause_prev[177] & ~x[2] & ~x[8] & ~x[32] & ~x[37] & ~x[58];
			partial_clause[178] 	= partial_clause_prev[178] & ~x[12];
			partial_clause[179] 	= partial_clause_prev[179] & ~x[10] & ~x[53];
			partial_clause[180] 	= partial_clause_prev[180] & ~x[34];
			partial_clause[181] 	= partial_clause_prev[181] & 1'b1;
			partial_clause[182] 	= partial_clause_prev[182] & ~x[23] & ~x[41] & ~x[50];
			partial_clause[183] 	= partial_clause_prev[183] & ~x[4] & ~x[5] & ~x[15] & ~x[16] & ~x[31] & ~x[36] & ~x[38] & ~x[42] & ~x[44] & ~x[45] & ~x[62];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[4] & ~x[11] & ~x[15] & ~x[31] & ~x[39] & ~x[43] & ~x[44] & ~x[62];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[33] & ~x[45];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[5] & ~x[6] & ~x[17] & ~x[39] & ~x[60] & ~x[63];
			partial_clause[187] 	= partial_clause_prev[187] & ~x[14] & ~x[19] & ~x[37] & ~x[39] & ~x[41] & ~x[50] & ~x[51];
			partial_clause[188] 	= partial_clause_prev[188] & x[30] & x[53];
			partial_clause[189] 	= partial_clause_prev[189] & 1'b1;
			partial_clause[190] 	= partial_clause_prev[190] & ~x[35] & ~x[40] & ~x[58];
			partial_clause[191] 	= partial_clause_prev[191] & ~x[12];
			partial_clause[192] 	= partial_clause_prev[192] & ~x[17] & ~x[45] & ~x[46];
			partial_clause[193] 	= partial_clause_prev[193] & ~x[6] & ~x[14] & ~x[40] & ~x[62];
			partial_clause[194] 	= partial_clause_prev[194] & ~x[39];
			partial_clause[195] 	= partial_clause_prev[195] & ~x[2] & ~x[10] & ~x[19] & ~x[35] & ~x[39] & ~x[45] & ~x[56] & ~x[57] & ~x[58] & ~x[63];
			partial_clause[196] 	= partial_clause_prev[196] & ~x[28] & ~x[47];
			partial_clause[197] 	= partial_clause_prev[197] & ~x[6] & ~x[7] & ~x[9] & ~x[13] & ~x[18] & ~x[39] & ~x[40] & ~x[42] & ~x[43] & ~x[44] & ~x[46];
			partial_clause[198] 	= partial_clause_prev[198] & ~x[30] & ~x[31];
			partial_clause[199] 	= partial_clause_prev[199] & 1'b1;
			partial_clause[200] 	= partial_clause_prev[200] & ~x[13] & ~x[39];
			partial_clause[201] 	= partial_clause_prev[201] & ~x[0] & ~x[30] & ~x[36] & ~x[41] & ~x[57] & ~x[58];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[9] & ~x[10] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[36] & ~x[38] & ~x[41] & ~x[62];
			partial_clause[203] 	= partial_clause_prev[203] & ~x[4] & ~x[34];
			partial_clause[204] 	= partial_clause_prev[204] & ~x[13] & ~x[15] & ~x[16] & ~x[17] & ~x[21] & ~x[33] & ~x[42] & ~x[46];
			partial_clause[205] 	= partial_clause_prev[205] & ~x[57] & ~x[62];
			partial_clause[206] 	= partial_clause_prev[206] & ~x[9] & ~x[14] & ~x[35] & ~x[36] & ~x[39] & ~x[63];
			partial_clause[207] 	= partial_clause_prev[207] & ~x[3] & ~x[8] & ~x[47] & ~x[49] & ~x[61] & ~x[63];
			partial_clause[208] 	= partial_clause_prev[208] & ~x[5] & ~x[38];
			partial_clause[209] 	= partial_clause_prev[209] & ~x[3] & ~x[57];
			partial_clause[210] 	= partial_clause_prev[210] & ~x[7] & ~x[9] & ~x[35] & ~x[61];
			partial_clause[211] 	= partial_clause_prev[211] & 1'b1;
			partial_clause[212] 	= partial_clause_prev[212] & ~x[5] & ~x[12] & ~x[14] & ~x[43];
			partial_clause[213] 	= partial_clause_prev[213] & ~x[4] & x[47] & ~x[58];
			partial_clause[214] 	= partial_clause_prev[214] & 1'b1;
			partial_clause[215] 	= partial_clause_prev[215] & 1'b1;
			partial_clause[216] 	= partial_clause_prev[216] & 1'b1;
			partial_clause[217] 	= partial_clause_prev[217] & ~x[41] & ~x[42] & ~x[44] & ~x[47];
			partial_clause[218] 	= partial_clause_prev[218] & ~x[7];
			partial_clause[219] 	= partial_clause_prev[219] & ~x[47] & ~x[49];
			partial_clause[220] 	= partial_clause_prev[220] & ~x[7] & ~x[9] & ~x[11] & ~x[13] & ~x[14] & ~x[15] & ~x[17] & ~x[32] & ~x[37] & ~x[38] & ~x[40] & ~x[43];
			partial_clause[221] 	= partial_clause_prev[221] & ~x[9] & ~x[15] & ~x[19] & ~x[40] & ~x[46];
			partial_clause[222] 	= partial_clause_prev[222] & 1'b1;
			partial_clause[223] 	= partial_clause_prev[223] & ~x[15] & ~x[28] & ~x[29] & ~x[32] & ~x[36];
			partial_clause[224] 	= partial_clause_prev[224] & ~x[7] & ~x[13] & ~x[34] & ~x[35] & ~x[46] & ~x[61];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[41];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[10] & ~x[16] & ~x[21] & ~x[23] & ~x[24] & ~x[38] & ~x[39] & ~x[41] & ~x[43] & ~x[44] & ~x[45] & ~x[48] & ~x[50] & ~x[52];
			partial_clause[227] 	= partial_clause_prev[227] & ~x[10] & ~x[51];
			partial_clause[228] 	= partial_clause_prev[228] & ~x[5] & ~x[10] & ~x[11] & ~x[16] & ~x[32] & ~x[36] & ~x[39];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[15] & ~x[36] & ~x[40] & ~x[41] & x[52] & x[53] & ~x[59] & ~x[63];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[8] & ~x[10] & ~x[12] & ~x[15] & ~x[33] & ~x[34] & ~x[35] & ~x[37] & ~x[39] & ~x[40] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[231] 	= partial_clause_prev[231] & ~x[7] & ~x[8] & ~x[10] & ~x[14] & ~x[36];
			partial_clause[232] 	= partial_clause_prev[232] & 1'b1;
			partial_clause[233] 	= partial_clause_prev[233] & 1'b1;
			partial_clause[234] 	= partial_clause_prev[234] & ~x[56];
			partial_clause[235] 	= partial_clause_prev[235] & 1'b1;
			partial_clause[236] 	= partial_clause_prev[236] & 1'b1;
			partial_clause[237] 	= partial_clause_prev[237] & 1'b1;
			partial_clause[238] 	= partial_clause_prev[238] & 1'b1;
			partial_clause[239] 	= partial_clause_prev[239] & ~x[10] & ~x[12];
			partial_clause[240] 	= partial_clause_prev[240] & ~x[3] & ~x[9] & ~x[46];
			partial_clause[241] 	= partial_clause_prev[241] & ~x[8] & ~x[14] & ~x[21] & ~x[23] & ~x[25] & ~x[44] & ~x[49];
			partial_clause[242] 	= partial_clause_prev[242] & ~x[8] & ~x[42] & ~x[43] & ~x[59] & ~x[62];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[10] & ~x[11] & ~x[14];
			partial_clause[244] 	= partial_clause_prev[244] & ~x[21] & ~x[22];
			partial_clause[245] 	= partial_clause_prev[245] & 1'b1;
			partial_clause[246] 	= partial_clause_prev[246] & ~x[10] & ~x[16];
			partial_clause[247] 	= partial_clause_prev[247] & ~x[4] & ~x[6] & ~x[8] & ~x[12] & ~x[13] & ~x[14] & ~x[16] & ~x[17] & ~x[34] & ~x[39] & ~x[40] & ~x[42] & ~x[45] & ~x[58] & ~x[60];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[18] & ~x[19] & ~x[33] & ~x[34] & ~x[37] & ~x[38] & ~x[43] & ~x[62] & ~x[63];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[38] & ~x[39];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[3] & ~x[4] & ~x[6] & ~x[8] & ~x[9] & ~x[11] & ~x[12] & ~x[14] & ~x[15] & ~x[17] & ~x[30] & ~x[31] & ~x[32] & ~x[35] & ~x[36] & ~x[38] & ~x[41] & ~x[42] & ~x[46] & ~x[58] & ~x[60];
			partial_clause[251] 	= partial_clause_prev[251] & ~x[0] & ~x[40];
			partial_clause[252] 	= partial_clause_prev[252] & ~x[8] & ~x[13] & ~x[16] & ~x[19] & ~x[36] & ~x[37] & ~x[38] & ~x[40] & ~x[45] & ~x[46] & ~x[47];
			partial_clause[253] 	= partial_clause_prev[253] & 1'b1;
			partial_clause[254] 	= partial_clause_prev[254] & ~x[18] & ~x[45];
			partial_clause[255] 	= partial_clause_prev[255] & ~x[14] & ~x[44];
			partial_clause[256] 	= partial_clause_prev[256] & 1'b1;
			partial_clause[257] 	= partial_clause_prev[257] & ~x[34];
			partial_clause[258] 	= partial_clause_prev[258] & ~x[6] & ~x[8] & ~x[18] & ~x[40] & ~x[47];
			partial_clause[259] 	= partial_clause_prev[259] & 1'b1;
			partial_clause[260] 	= partial_clause_prev[260] & ~x[10] & ~x[13] & ~x[15] & ~x[42];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[8] & ~x[11] & ~x[31] & ~x[33] & ~x[41];
			partial_clause[262] 	= partial_clause_prev[262] & ~x[10] & ~x[47] & x[55];
			partial_clause[263] 	= partial_clause_prev[263] & ~x[1] & ~x[20] & ~x[35];
			partial_clause[264] 	= partial_clause_prev[264] & ~x[2] & ~x[7] & ~x[10] & ~x[15] & ~x[35] & ~x[58];
			partial_clause[265] 	= partial_clause_prev[265] & x[24];
			partial_clause[266] 	= partial_clause_prev[266] & ~x[10] & ~x[11] & ~x[12] & ~x[32] & ~x[45] & ~x[59] & ~x[62];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[9] & ~x[10] & ~x[14] & ~x[15] & ~x[16] & ~x[35] & ~x[46] & ~x[47] & ~x[59] & ~x[60];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[9] & ~x[13] & ~x[15] & ~x[38] & ~x[39] & ~x[40];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[8] & ~x[10] & ~x[12] & ~x[13] & ~x[34] & ~x[35] & ~x[37] & ~x[38] & ~x[39] & ~x[43] & ~x[59] & ~x[60] & ~x[62];
			partial_clause[270] 	= partial_clause_prev[270] & 1'b1;
			partial_clause[271] 	= partial_clause_prev[271] & ~x[46];
			partial_clause[272] 	= partial_clause_prev[272] & ~x[7] & ~x[10] & ~x[12] & ~x[14] & ~x[15] & ~x[63];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[7] & ~x[8] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[17] & ~x[18] & ~x[20] & ~x[35] & ~x[39] & ~x[40] & ~x[43] & ~x[47] & ~x[49];
			partial_clause[274] 	= partial_clause_prev[274] & ~x[9] & ~x[12];
			partial_clause[275] 	= partial_clause_prev[275] & ~x[9];
			partial_clause[276] 	= partial_clause_prev[276] & ~x[14] & ~x[19] & ~x[43];
			partial_clause[277] 	= partial_clause_prev[277] & ~x[33] & ~x[39];
			partial_clause[278] 	= partial_clause_prev[278] & 1'b1;
			partial_clause[279] 	= partial_clause_prev[279] & ~x[3] & ~x[4] & ~x[7] & ~x[8] & ~x[11] & ~x[12] & ~x[13] & ~x[17] & ~x[19] & ~x[31] & ~x[34] & ~x[36] & ~x[37] & ~x[38] & ~x[39] & ~x[43] & ~x[44] & ~x[46] & ~x[47];
			partial_clause[280] 	= partial_clause_prev[280] & 1'b1;
			partial_clause[281] 	= partial_clause_prev[281] & ~x[13] & ~x[16] & ~x[45] & ~x[62];
			partial_clause[282] 	= partial_clause_prev[282] & ~x[12] & ~x[15] & ~x[16] & ~x[17] & x[50];
			partial_clause[283] 	= partial_clause_prev[283] & ~x[56];
			partial_clause[284] 	= partial_clause_prev[284] & 1'b1;
			partial_clause[285] 	= partial_clause_prev[285] & 1'b1;
			partial_clause[286] 	= partial_clause_prev[286] & ~x[2] & ~x[27] & ~x[55];
			partial_clause[287] 	= partial_clause_prev[287] & ~x[6] & ~x[8] & ~x[13] & ~x[15] & ~x[33] & ~x[35] & ~x[36] & ~x[37] & ~x[41] & ~x[44] & ~x[60];
			partial_clause[288] 	= partial_clause_prev[288] & ~x[6];
			partial_clause[289] 	= partial_clause_prev[289] & ~x[42];
			partial_clause[290] 	= partial_clause_prev[290] & 1'b1;
			partial_clause[291] 	= partial_clause_prev[291] & 1'b1;
			partial_clause[292] 	= partial_clause_prev[292] & ~x[1] & ~x[7] & ~x[8] & ~x[18] & ~x[30] & ~x[41] & ~x[46];
			partial_clause[293] 	= partial_clause_prev[293] & ~x[4] & ~x[5] & ~x[10] & ~x[16] & ~x[18] & ~x[43];
			partial_clause[294] 	= partial_clause_prev[294] & 1'b1;
			partial_clause[295] 	= partial_clause_prev[295] & ~x[9] & ~x[14];
			partial_clause[296] 	= partial_clause_prev[296] & ~x[15];
			partial_clause[297] 	= partial_clause_prev[297] & ~x[8] & ~x[16] & ~x[18] & ~x[27];
			partial_clause[298] 	= partial_clause_prev[298] & 1'b1;
			partial_clause[299] 	= partial_clause_prev[299] & ~x[6] & ~x[7] & ~x[14] & ~x[15] & ~x[62];
			partial_clause[300] 	= partial_clause_prev[300] & 1'b1;
			partial_clause[301] 	= partial_clause_prev[301] & ~x[3] & ~x[19] & ~x[20] & ~x[32] & ~x[62];
			partial_clause[302] 	= partial_clause_prev[302] & ~x[11];
			partial_clause[303] 	= partial_clause_prev[303] & ~x[4] & ~x[19] & ~x[45];
			partial_clause[304] 	= partial_clause_prev[304] & ~x[44];
			partial_clause[305] 	= partial_clause_prev[305] & ~x[15] & ~x[33] & ~x[37] & ~x[63];
			partial_clause[306] 	= partial_clause_prev[306] & ~x[13] & ~x[16] & ~x[21] & ~x[32] & ~x[33] & ~x[39] & ~x[41] & ~x[45] & ~x[47] & ~x[48] & ~x[50] & ~x[58] & ~x[60] & ~x[61];
			partial_clause[307] 	= partial_clause_prev[307] & ~x[3] & ~x[12] & ~x[40] & ~x[44] & ~x[55];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[7] & ~x[8] & ~x[13] & ~x[38] & ~x[49] & ~x[63];
			partial_clause[309] 	= partial_clause_prev[309] & ~x[15];
			partial_clause[310] 	= partial_clause_prev[310] & 1'b1;
			partial_clause[311] 	= partial_clause_prev[311] & ~x[17] & ~x[27] & ~x[54];
			partial_clause[312] 	= partial_clause_prev[312] & ~x[32] & ~x[41] & ~x[60];
			partial_clause[313] 	= partial_clause_prev[313] & ~x[52];
			partial_clause[314] 	= partial_clause_prev[314] & 1'b1;
			partial_clause[315] 	= partial_clause_prev[315] & ~x[17] & ~x[41] & ~x[42];
			partial_clause[316] 	= partial_clause_prev[316] & ~x[13] & ~x[14] & ~x[16] & ~x[35] & ~x[36] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[46] & ~x[47] & ~x[62];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[10] & ~x[19];
			partial_clause[318] 	= partial_clause_prev[318] & ~x[4] & ~x[13] & ~x[15] & ~x[62];
			partial_clause[319] 	= partial_clause_prev[319] & ~x[9] & ~x[12] & ~x[38];
			partial_clause[320] 	= partial_clause_prev[320] & ~x[15] & ~x[62];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[5] & ~x[13] & ~x[15] & ~x[35];
			partial_clause[322] 	= partial_clause_prev[322] & ~x[4] & ~x[37] & ~x[62];
			partial_clause[323] 	= partial_clause_prev[323] & ~x[34] & ~x[42] & ~x[44] & ~x[46];
			partial_clause[324] 	= partial_clause_prev[324] & ~x[15] & ~x[16];
			partial_clause[325] 	= partial_clause_prev[325] & ~x[3] & ~x[5] & ~x[6] & ~x[8] & ~x[11] & ~x[13] & x[27] & ~x[31] & ~x[33] & ~x[34] & ~x[43] & ~x[59] & ~x[60];
			partial_clause[326] 	= partial_clause_prev[326] & ~x[12] & ~x[37];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[34] & ~x[49] & ~x[59];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[62] & ~x[63];
			partial_clause[329] 	= partial_clause_prev[329] & 1'b1;
			partial_clause[330] 	= partial_clause_prev[330] & ~x[15] & x[52];
			partial_clause[331] 	= partial_clause_prev[331] & ~x[59];
			partial_clause[332] 	= partial_clause_prev[332] & ~x[12] & ~x[44] & ~x[62];
			partial_clause[333] 	= partial_clause_prev[333] & ~x[63];
			partial_clause[334] 	= partial_clause_prev[334] & ~x[9] & x[29];
			partial_clause[335] 	= partial_clause_prev[335] & ~x[8];
			partial_clause[336] 	= partial_clause_prev[336] & 1'b1;
			partial_clause[337] 	= partial_clause_prev[337] & ~x[11] & ~x[12] & ~x[14] & ~x[41] & ~x[43];
			partial_clause[338] 	= partial_clause_prev[338] & x[0];
			partial_clause[339] 	= partial_clause_prev[339] & ~x[6] & ~x[11] & ~x[37] & ~x[38] & ~x[59] & ~x[62];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[15] & ~x[16] & ~x[18] & ~x[35] & ~x[46] & ~x[48];
			partial_clause[341] 	= partial_clause_prev[341] & 1'b1;
			partial_clause[342] 	= partial_clause_prev[342] & ~x[36] & ~x[63];
			partial_clause[343] 	= partial_clause_prev[343] & ~x[35] & ~x[41] & ~x[62];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[5] & ~x[15] & ~x[44];
			partial_clause[345] 	= partial_clause_prev[345] & 1'b1;
			partial_clause[346] 	= partial_clause_prev[346] & 1'b1;
			partial_clause[347] 	= partial_clause_prev[347] & ~x[14];
			partial_clause[348] 	= partial_clause_prev[348] & x[32];
			partial_clause[349] 	= partial_clause_prev[349] & ~x[8] & ~x[11];
			partial_clause[350] 	= partial_clause_prev[350] & ~x[9] & ~x[12] & ~x[15] & ~x[16] & ~x[18] & ~x[34] & ~x[37] & ~x[40] & ~x[41] & ~x[44] & ~x[45] & ~x[47] & ~x[49] & ~x[63];
			partial_clause[351] 	= partial_clause_prev[351] & 1'b1;
			partial_clause[352] 	= partial_clause_prev[352] & 1'b1;
			partial_clause[353] 	= partial_clause_prev[353] & 1'b1;
			partial_clause[354] 	= partial_clause_prev[354] & 1'b1;
			partial_clause[355] 	= partial_clause_prev[355] & ~x[7] & ~x[9] & ~x[16] & ~x[61];
			partial_clause[356] 	= partial_clause_prev[356] & ~x[35] & ~x[41];
			partial_clause[357] 	= partial_clause_prev[357] & ~x[62];
			partial_clause[358] 	= partial_clause_prev[358] & ~x[13] & ~x[14] & ~x[20] & ~x[22] & ~x[37] & ~x[49] & ~x[50] & ~x[61];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[16] & ~x[20] & ~x[41];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[13] & ~x[15] & ~x[18] & ~x[21] & ~x[22] & ~x[34] & ~x[40] & ~x[43] & ~x[44] & ~x[45] & ~x[49];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[13] & ~x[16] & ~x[40] & ~x[41] & ~x[45] & ~x[61];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[0] & ~x[13] & ~x[39] & ~x[57];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[14] & ~x[40] & ~x[45] & ~x[49];
			partial_clause[364] 	= partial_clause_prev[364] & ~x[6] & ~x[13] & x[24] & ~x[31] & ~x[35];
			partial_clause[365] 	= partial_clause_prev[365] & 1'b1;
			partial_clause[366] 	= partial_clause_prev[366] & ~x[9] & ~x[10] & ~x[14] & ~x[17] & ~x[18] & ~x[41] & ~x[43];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[13] & ~x[39];
			partial_clause[368] 	= partial_clause_prev[368] & 1'b1;
			partial_clause[369] 	= partial_clause_prev[369] & ~x[16] & ~x[37] & ~x[46];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[2] & ~x[12] & ~x[20] & ~x[29] & ~x[57] & ~x[61];
			partial_clause[371] 	= partial_clause_prev[371] & ~x[6] & ~x[45];
			partial_clause[372] 	= partial_clause_prev[372] & ~x[3] & ~x[7] & ~x[33] & ~x[34] & ~x[43];
			partial_clause[373] 	= partial_clause_prev[373] & ~x[46];
			partial_clause[374] 	= partial_clause_prev[374] & ~x[42];
			partial_clause[375] 	= partial_clause_prev[375] & ~x[7] & ~x[34];
			partial_clause[376] 	= partial_clause_prev[376] & ~x[7] & ~x[19] & ~x[20] & ~x[44] & ~x[45];
			partial_clause[377] 	= partial_clause_prev[377] & x[21] & ~x[40];
			partial_clause[378] 	= partial_clause_prev[378] & ~x[11];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[41] & ~x[63];
			partial_clause[380] 	= partial_clause_prev[380] & ~x[19];
			partial_clause[381] 	= partial_clause_prev[381] & ~x[12] & ~x[35] & ~x[38] & ~x[39];
			partial_clause[382] 	= partial_clause_prev[382] & 1'b1;
			partial_clause[383] 	= partial_clause_prev[383] & ~x[3] & ~x[31];
			partial_clause[384] 	= partial_clause_prev[384] & 1'b1;
			partial_clause[385] 	= partial_clause_prev[385] & 1'b1;
			partial_clause[386] 	= partial_clause_prev[386] & x[23];
			partial_clause[387] 	= partial_clause_prev[387] & ~x[12] & ~x[16] & ~x[17] & ~x[38] & ~x[40] & ~x[41] & ~x[42] & ~x[44];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[10] & ~x[15] & ~x[38] & ~x[39] & ~x[42] & ~x[43];
			partial_clause[389] 	= partial_clause_prev[389] & 1'b1;
			partial_clause[390] 	= partial_clause_prev[390] & ~x[5] & ~x[6] & ~x[8] & ~x[12] & ~x[38] & ~x[41] & ~x[61] & ~x[62];
			partial_clause[391] 	= partial_clause_prev[391] & 1'b1;
			partial_clause[392] 	= partial_clause_prev[392] & 1'b1;
			partial_clause[393] 	= partial_clause_prev[393] & 1'b1;
			partial_clause[394] 	= partial_clause_prev[394] & ~x[38];
			partial_clause[395] 	= partial_clause_prev[395] & x[26] & ~x[61] & ~x[62];
			partial_clause[396] 	= partial_clause_prev[396] & ~x[58] & ~x[60];
			partial_clause[397] 	= partial_clause_prev[397] & 1'b1;
			partial_clause[398] 	= partial_clause_prev[398] & 1'b1;
			partial_clause[399] 	= partial_clause_prev[399] & 1'b1;
			partial_clause[400] 	= partial_clause_prev[400] & ~x[7] & ~x[9] & ~x[11] & ~x[16] & ~x[19] & ~x[45] & ~x[47] & ~x[62];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[5] & ~x[8] & ~x[13] & ~x[34] & ~x[38] & ~x[39] & ~x[41] & ~x[44] & ~x[45] & ~x[59] & ~x[63];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[9] & ~x[12] & ~x[17] & ~x[35] & ~x[44];
			partial_clause[403] 	= partial_clause_prev[403] & ~x[9] & ~x[12] & ~x[19] & ~x[40] & ~x[46] & ~x[49];
			partial_clause[404] 	= partial_clause_prev[404] & 1'b1;
			partial_clause[405] 	= partial_clause_prev[405] & ~x[14] & ~x[42] & ~x[61];
			partial_clause[406] 	= partial_clause_prev[406] & ~x[33] & ~x[41];
			partial_clause[407] 	= partial_clause_prev[407] & 1'b1;
			partial_clause[408] 	= partial_clause_prev[408] & 1'b1;
			partial_clause[409] 	= partial_clause_prev[409] & ~x[4] & ~x[5] & ~x[12] & ~x[13] & ~x[15] & ~x[31] & ~x[46] & ~x[58] & ~x[62];
			partial_clause[410] 	= partial_clause_prev[410] & ~x[6] & ~x[34] & ~x[43];
			partial_clause[411] 	= partial_clause_prev[411] & ~x[12] & ~x[52];
			partial_clause[412] 	= partial_clause_prev[412] & ~x[5] & ~x[8] & ~x[11] & ~x[15] & ~x[36] & ~x[41] & ~x[42] & ~x[45];
			partial_clause[413] 	= partial_clause_prev[413] & x[52];
			partial_clause[414] 	= partial_clause_prev[414] & ~x[5] & ~x[10] & ~x[14] & ~x[16] & ~x[37] & ~x[39];
			partial_clause[415] 	= partial_clause_prev[415] & ~x[19] & ~x[44] & ~x[45];
			partial_clause[416] 	= partial_clause_prev[416] & ~x[3] & ~x[13] & ~x[15] & x[23] & ~x[32] & ~x[42] & ~x[43] & ~x[58] & ~x[59];
			partial_clause[417] 	= partial_clause_prev[417] & ~x[8] & ~x[37] & ~x[61];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[5] & ~x[7] & ~x[13] & ~x[18] & ~x[19] & ~x[21] & ~x[32] & ~x[35] & ~x[36] & ~x[40] & ~x[42] & ~x[43] & ~x[45];
			partial_clause[419] 	= partial_clause_prev[419] & 1'b1;
			partial_clause[420] 	= partial_clause_prev[420] & 1'b1;
			partial_clause[421] 	= partial_clause_prev[421] & ~x[8] & ~x[9] & ~x[11] & ~x[16] & ~x[17] & ~x[37] & ~x[39] & ~x[41] & ~x[42] & ~x[44] & ~x[45] & ~x[46];
			partial_clause[422] 	= partial_clause_prev[422] & ~x[7] & ~x[13] & ~x[20] & ~x[38];
			partial_clause[423] 	= partial_clause_prev[423] & ~x[38];
			partial_clause[424] 	= partial_clause_prev[424] & ~x[10];
			partial_clause[425] 	= partial_clause_prev[425] & 1'b1;
			partial_clause[426] 	= partial_clause_prev[426] & ~x[9] & ~x[11] & ~x[13] & ~x[36] & ~x[37] & ~x[40] & ~x[45] & ~x[62];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[12];
			partial_clause[428] 	= partial_clause_prev[428] & ~x[13] & ~x[44] & ~x[51] & ~x[52] & ~x[55] & ~x[56] & ~x[57] & ~x[63];
			partial_clause[429] 	= partial_clause_prev[429] & 1'b1;
			partial_clause[430] 	= partial_clause_prev[430] & ~x[4] & ~x[17] & ~x[32] & ~x[35] & ~x[38] & ~x[39] & ~x[41] & ~x[42] & ~x[43];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[9] & ~x[10];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[8] & ~x[41] & ~x[62] & ~x[63];
			partial_clause[433] 	= partial_clause_prev[433] & ~x[39];
			partial_clause[434] 	= partial_clause_prev[434] & ~x[18] & ~x[23];
			partial_clause[435] 	= partial_clause_prev[435] & ~x[8] & ~x[11] & ~x[32] & ~x[35] & ~x[36] & ~x[37] & ~x[42] & ~x[44];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[40] & ~x[41];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[7] & ~x[15] & ~x[31] & ~x[32] & ~x[44] & ~x[60] & ~x[63];
			partial_clause[438] 	= partial_clause_prev[438] & ~x[17] & ~x[41];
			partial_clause[439] 	= partial_clause_prev[439] & ~x[63];
			partial_clause[440] 	= partial_clause_prev[440] & x[24];
			partial_clause[441] 	= partial_clause_prev[441] & ~x[13];
			partial_clause[442] 	= partial_clause_prev[442] & 1'b1;
			partial_clause[443] 	= partial_clause_prev[443] & ~x[6] & ~x[34] & ~x[44];
			partial_clause[444] 	= partial_clause_prev[444] & 1'b1;
			partial_clause[445] 	= partial_clause_prev[445] & 1'b1;
			partial_clause[446] 	= partial_clause_prev[446] & ~x[10] & ~x[63];
			partial_clause[447] 	= partial_clause_prev[447] & ~x[8] & ~x[11] & ~x[12] & ~x[37] & ~x[38] & ~x[39] & ~x[41] & x[55];
			partial_clause[448] 	= partial_clause_prev[448] & 1'b1;
			partial_clause[449] 	= partial_clause_prev[449] & ~x[13] & ~x[38];
			partial_clause[450] 	= partial_clause_prev[450] & ~x[3] & ~x[7] & ~x[8] & ~x[12] & ~x[34] & ~x[46];
			partial_clause[451] 	= partial_clause_prev[451] & 1'b1;
			partial_clause[452] 	= partial_clause_prev[452] & 1'b1;
			partial_clause[453] 	= partial_clause_prev[453] & ~x[10] & ~x[24] & ~x[33];
			partial_clause[454] 	= partial_clause_prev[454] & 1'b1;
			partial_clause[455] 	= partial_clause_prev[455] & ~x[8] & ~x[9] & ~x[17] & ~x[19] & ~x[33];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[13] & ~x[35] & ~x[41] & ~x[43] & ~x[44] & x[52] & x[53] & ~x[59] & ~x[62] & ~x[63];
			partial_clause[457] 	= partial_clause_prev[457] & ~x[15];
			partial_clause[458] 	= partial_clause_prev[458] & ~x[8] & ~x[38] & ~x[61] & ~x[62];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[9] & ~x[30] & ~x[39] & ~x[57] & ~x[58];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[13] & ~x[15] & ~x[32] & ~x[34] & ~x[37] & ~x[39] & ~x[60];
			partial_clause[461] 	= partial_clause_prev[461] & ~x[24] & ~x[37] & ~x[38] & ~x[41];
			partial_clause[462] 	= partial_clause_prev[462] & ~x[10] & ~x[40];
			partial_clause[463] 	= partial_clause_prev[463] & 1'b1;
			partial_clause[464] 	= partial_clause_prev[464] & ~x[38] & ~x[39] & ~x[40] & ~x[61];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[10] & ~x[11] & ~x[40] & ~x[41];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[12] & ~x[15] & ~x[39] & ~x[43];
			partial_clause[467] 	= partial_clause_prev[467] & 1'b1;
			partial_clause[468] 	= partial_clause_prev[468] & ~x[5] & ~x[8] & ~x[32] & ~x[35] & ~x[60];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[8];
			partial_clause[470] 	= partial_clause_prev[470] & 1'b1;
			partial_clause[471] 	= partial_clause_prev[471] & ~x[3] & ~x[4] & ~x[12] & ~x[31] & ~x[33] & ~x[45] & ~x[57] & ~x[58] & ~x[59] & ~x[60] & ~x[63];
			partial_clause[472] 	= partial_clause_prev[472] & ~x[16] & ~x[31] & ~x[44] & ~x[58] & ~x[63];
			partial_clause[473] 	= partial_clause_prev[473] & ~x[9] & ~x[34] & ~x[39] & ~x[41];
			partial_clause[474] 	= partial_clause_prev[474] & ~x[26] & ~x[27];
			partial_clause[475] 	= partial_clause_prev[475] & ~x[16] & ~x[41];
			partial_clause[476] 	= partial_clause_prev[476] & x[25] & ~x[52];
			partial_clause[477] 	= partial_clause_prev[477] & ~x[42];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[12] & ~x[19] & ~x[36] & ~x[46] & ~x[63];
			partial_clause[479] 	= partial_clause_prev[479] & 1'b1;
			partial_clause[480] 	= partial_clause_prev[480] & ~x[7] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[17] & ~x[33] & ~x[34] & ~x[37] & ~x[38] & ~x[39] & ~x[41] & ~x[42] & ~x[43] & ~x[45] & ~x[63];
			partial_clause[481] 	= partial_clause_prev[481] & 1'b1;
			partial_clause[482] 	= partial_clause_prev[482] & ~x[9] & ~x[40] & ~x[46];
			partial_clause[483] 	= partial_clause_prev[483] & ~x[4] & ~x[9];
			partial_clause[484] 	= partial_clause_prev[484] & ~x[42];
			partial_clause[485] 	= partial_clause_prev[485] & x[1] & ~x[35] & ~x[62];
			partial_clause[486] 	= partial_clause_prev[486] & ~x[10] & ~x[41];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[8] & ~x[16] & ~x[44] & ~x[63];
			partial_clause[488] 	= partial_clause_prev[488] & 1'b1;
			partial_clause[489] 	= partial_clause_prev[489] & ~x[53] & ~x[54];
			partial_clause[490] 	= partial_clause_prev[490] & 1'b1;
			partial_clause[491] 	= partial_clause_prev[491] & 1'b1;
			partial_clause[492] 	= partial_clause_prev[492] & ~x[55];
			partial_clause[493] 	= partial_clause_prev[493] & 1'b1;
			partial_clause[494] 	= partial_clause_prev[494] & ~x[9] & ~x[12] & ~x[39] & x[52] & ~x[62];
			partial_clause[495] 	= partial_clause_prev[495] & ~x[11] & ~x[12] & ~x[15] & ~x[39];
			partial_clause[496] 	= partial_clause_prev[496] & ~x[51];
			partial_clause[497] 	= partial_clause_prev[497] & ~x[20];
			partial_clause[498] 	= partial_clause_prev[498] & x[49];
			partial_clause[499] 	= partial_clause_prev[499] & ~x[12];
		end
	end
endmodule


module HCB_10 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[0] & ~x[3] & ~x[4] & ~x[5] & ~x[29] & ~x[30] & ~x[31] & ~x[56] & ~x[57] & ~x[61] & ~x[62];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[1] & ~x[2] & ~x[8] & ~x[22] & ~x[35] & ~x[36] & ~x[40];
			partial_clause[2] 	= partial_clause_prev[2] & ~x[27];
			partial_clause[3] 	= partial_clause_prev[3] & ~x[28] & ~x[51] & ~x[52];
			partial_clause[4] 	= partial_clause_prev[4] & 1'b1;
			partial_clause[5] 	= partial_clause_prev[5] & ~x[5] & ~x[10] & ~x[11] & ~x[28] & ~x[30] & ~x[32] & ~x[33] & ~x[35];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[1] & ~x[27] & ~x[42] & ~x[50] & ~x[51] & ~x[60];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[4] & ~x[9] & ~x[11] & ~x[40] & ~x[55] & ~x[58] & ~x[63];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[5] & ~x[20] & ~x[23] & ~x[26] & ~x[29] & ~x[30] & ~x[34] & ~x[60];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[1] & ~x[4] & ~x[8] & ~x[11] & ~x[26] & ~x[29] & ~x[34] & ~x[36] & ~x[52] & ~x[57] & ~x[59];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[3] & ~x[22] & ~x[25] & ~x[27] & ~x[29] & ~x[58] & ~x[59];
			partial_clause[11] 	= partial_clause_prev[11] & ~x[2] & ~x[4] & ~x[20] & ~x[22] & ~x[30] & ~x[32] & ~x[49] & ~x[50] & ~x[52] & ~x[59] & ~x[63];
			partial_clause[12] 	= partial_clause_prev[12] & ~x[8] & ~x[34] & ~x[35] & ~x[37];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[0] & ~x[7] & ~x[8] & ~x[22] & ~x[23] & ~x[26] & ~x[32] & ~x[33] & ~x[50] & ~x[54] & ~x[59] & ~x[60] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[14] 	= partial_clause_prev[14] & 1'b1;
			partial_clause[15] 	= partial_clause_prev[15] & ~x[14] & ~x[16];
			partial_clause[16] 	= partial_clause_prev[16] & ~x[25] & ~x[34] & ~x[35] & ~x[62];
			partial_clause[17] 	= partial_clause_prev[17] & ~x[4] & x[18] & ~x[32];
			partial_clause[18] 	= partial_clause_prev[18] & ~x[1] & ~x[28] & ~x[44] & ~x[49] & ~x[53] & ~x[56];
			partial_clause[19] 	= partial_clause_prev[19] & ~x[27] & ~x[30] & ~x[32] & ~x[34];
			partial_clause[20] 	= partial_clause_prev[20] & ~x[28] & ~x[43];
			partial_clause[21] 	= partial_clause_prev[21] & ~x[0] & ~x[33];
			partial_clause[22] 	= partial_clause_prev[22] & ~x[34] & ~x[38] & ~x[46] & ~x[48] & ~x[58];
			partial_clause[23] 	= partial_clause_prev[23] & ~x[1] & ~x[2] & ~x[4] & ~x[6] & ~x[9] & ~x[10] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & ~x[30] & ~x[31] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[38] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[45] & ~x[46] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[54] & ~x[56] & ~x[57] & ~x[60] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[3] & ~x[5] & ~x[6] & ~x[8] & ~x[10] & ~x[24] & ~x[26] & ~x[27] & ~x[28] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[35] & ~x[36] & ~x[37] & ~x[38] & ~x[40] & ~x[53] & ~x[54] & ~x[55] & ~x[57] & ~x[59] & ~x[61] & ~x[62];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[2] & ~x[3] & ~x[5] & ~x[6] & ~x[20] & ~x[22] & ~x[24] & ~x[25] & ~x[28] & ~x[30] & ~x[31] & ~x[32] & ~x[48] & ~x[50] & ~x[52] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[26] 	= partial_clause_prev[26] & 1'b1;
			partial_clause[27] 	= partial_clause_prev[27] & ~x[4] & ~x[8] & ~x[23] & ~x[32] & ~x[35] & ~x[36] & ~x[49] & ~x[50] & ~x[51] & ~x[54] & ~x[56] & ~x[60];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[8] & ~x[35] & ~x[60];
			partial_clause[29] 	= partial_clause_prev[29] & ~x[7] & ~x[28] & ~x[34];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[6] & ~x[7] & ~x[22] & ~x[25] & ~x[26] & ~x[52] & ~x[63];
			partial_clause[31] 	= partial_clause_prev[31] & ~x[35];
			partial_clause[32] 	= partial_clause_prev[32] & ~x[0] & ~x[1];
			partial_clause[33] 	= partial_clause_prev[33] & 1'b1;
			partial_clause[34] 	= partial_clause_prev[34] & ~x[1] & ~x[4] & ~x[6] & ~x[8] & ~x[10] & ~x[28] & ~x[31] & ~x[35] & ~x[37] & ~x[38] & ~x[54] & ~x[58] & ~x[60] & ~x[61] & ~x[63];
			partial_clause[35] 	= partial_clause_prev[35] & ~x[1] & ~x[30] & ~x[37];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[0] & ~x[2] & ~x[24] & ~x[28] & ~x[38] & ~x[41] & ~x[58] & ~x[59] & ~x[62];
			partial_clause[37] 	= partial_clause_prev[37] & ~x[36] & ~x[58];
			partial_clause[38] 	= partial_clause_prev[38] & ~x[3] & ~x[22] & ~x[34] & ~x[48] & ~x[50] & ~x[51] & ~x[52] & ~x[56] & ~x[63];
			partial_clause[39] 	= partial_clause_prev[39] & ~x[33] & ~x[42] & ~x[53];
			partial_clause[40] 	= partial_clause_prev[40] & ~x[6] & ~x[26];
			partial_clause[41] 	= partial_clause_prev[41] & 1'b1;
			partial_clause[42] 	= partial_clause_prev[42] & 1'b1;
			partial_clause[43] 	= partial_clause_prev[43] & ~x[1] & ~x[3] & ~x[10] & ~x[27] & ~x[56] & ~x[58] & ~x[63];
			partial_clause[44] 	= partial_clause_prev[44] & ~x[36] & ~x[57];
			partial_clause[45] 	= partial_clause_prev[45] & ~x[57];
			partial_clause[46] 	= partial_clause_prev[46] & ~x[0] & ~x[23] & ~x[26] & ~x[29] & ~x[50] & ~x[57];
			partial_clause[47] 	= partial_clause_prev[47] & ~x[23] & ~x[56];
			partial_clause[48] 	= partial_clause_prev[48] & 1'b1;
			partial_clause[49] 	= partial_clause_prev[49] & 1'b1;
			partial_clause[50] 	= partial_clause_prev[50] & ~x[55];
			partial_clause[51] 	= partial_clause_prev[51] & 1'b1;
			partial_clause[52] 	= partial_clause_prev[52] & ~x[36];
			partial_clause[53] 	= partial_clause_prev[53] & 1'b1;
			partial_clause[54] 	= partial_clause_prev[54] & ~x[4] & ~x[59];
			partial_clause[55] 	= partial_clause_prev[55] & ~x[45];
			partial_clause[56] 	= partial_clause_prev[56] & 1'b1;
			partial_clause[57] 	= partial_clause_prev[57] & ~x[4] & ~x[8] & ~x[22] & ~x[53] & ~x[58];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[7] & ~x[19] & ~x[32] & ~x[47] & ~x[49] & ~x[56];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[1] & ~x[12] & ~x[29] & ~x[31] & ~x[32] & ~x[36] & ~x[58] & ~x[60];
			partial_clause[60] 	= partial_clause_prev[60] & 1'b1;
			partial_clause[61] 	= partial_clause_prev[61] & ~x[4];
			partial_clause[62] 	= partial_clause_prev[62] & ~x[13] & ~x[14] & ~x[31] & ~x[35] & ~x[55];
			partial_clause[63] 	= partial_clause_prev[63] & ~x[1] & ~x[51];
			partial_clause[64] 	= partial_clause_prev[64] & 1'b1;
			partial_clause[65] 	= partial_clause_prev[65] & ~x[43];
			partial_clause[66] 	= partial_clause_prev[66] & 1'b1;
			partial_clause[67] 	= partial_clause_prev[67] & 1'b1;
			partial_clause[68] 	= partial_clause_prev[68] & ~x[9] & ~x[24] & ~x[27];
			partial_clause[69] 	= partial_clause_prev[69] & ~x[3] & ~x[7] & ~x[31] & ~x[32] & ~x[54] & ~x[55] & ~x[56];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[0] & ~x[2] & ~x[29] & ~x[35] & ~x[53];
			partial_clause[71] 	= partial_clause_prev[71] & ~x[61];
			partial_clause[72] 	= partial_clause_prev[72] & ~x[21];
			partial_clause[73] 	= partial_clause_prev[73] & ~x[28] & ~x[36];
			partial_clause[74] 	= partial_clause_prev[74] & ~x[1] & ~x[31] & ~x[33] & ~x[37] & ~x[55] & ~x[56];
			partial_clause[75] 	= partial_clause_prev[75] & ~x[50];
			partial_clause[76] 	= partial_clause_prev[76] & ~x[0] & ~x[8] & ~x[30] & ~x[31] & ~x[36] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[53];
			partial_clause[78] 	= partial_clause_prev[78] & ~x[52];
			partial_clause[79] 	= partial_clause_prev[79] & 1'b1;
			partial_clause[80] 	= partial_clause_prev[80] & 1'b1;
			partial_clause[81] 	= partial_clause_prev[81] & ~x[52] & ~x[60];
			partial_clause[82] 	= partial_clause_prev[82] & 1'b1;
			partial_clause[83] 	= partial_clause_prev[83] & 1'b1;
			partial_clause[84] 	= partial_clause_prev[84] & ~x[3] & ~x[7] & ~x[53] & ~x[61];
			partial_clause[85] 	= partial_clause_prev[85] & ~x[0] & ~x[4] & ~x[9] & ~x[30] & ~x[33] & ~x[53] & ~x[56] & ~x[60] & ~x[61] & ~x[63];
			partial_clause[86] 	= partial_clause_prev[86] & ~x[5] & ~x[6] & ~x[7] & ~x[26] & ~x[27] & ~x[50] & ~x[59] & ~x[60];
			partial_clause[87] 	= partial_clause_prev[87] & ~x[2] & ~x[8] & ~x[50] & ~x[53];
			partial_clause[88] 	= partial_clause_prev[88] & ~x[3] & ~x[4] & ~x[26] & ~x[34] & ~x[54];
			partial_clause[89] 	= partial_clause_prev[89] & ~x[4] & ~x[32] & ~x[34];
			partial_clause[90] 	= partial_clause_prev[90] & 1'b1;
			partial_clause[91] 	= partial_clause_prev[91] & ~x[25] & ~x[34];
			partial_clause[92] 	= partial_clause_prev[92] & ~x[3] & ~x[26] & ~x[57];
			partial_clause[93] 	= partial_clause_prev[93] & ~x[5] & ~x[10] & ~x[30] & ~x[32] & ~x[33] & ~x[34] & ~x[35] & ~x[37] & ~x[38] & ~x[41] & ~x[51] & ~x[54] & ~x[55] & ~x[56] & ~x[58] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[94] 	= partial_clause_prev[94] & 1'b1;
			partial_clause[95] 	= partial_clause_prev[95] & ~x[0] & ~x[2] & ~x[4] & ~x[35] & ~x[57] & ~x[61];
			partial_clause[96] 	= partial_clause_prev[96] & 1'b1;
			partial_clause[97] 	= partial_clause_prev[97] & ~x[3] & ~x[7] & ~x[10] & ~x[30] & ~x[31] & ~x[32] & ~x[38] & ~x[40] & ~x[55] & ~x[57] & ~x[58] & ~x[59] & ~x[61];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[0] & ~x[1] & ~x[9] & ~x[10] & ~x[12] & ~x[26] & ~x[32] & ~x[34] & ~x[36] & ~x[37] & ~x[40] & ~x[53] & ~x[58] & ~x[61];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[8] & ~x[9] & ~x[10] & ~x[11] & ~x[25] & ~x[26] & ~x[27] & ~x[28] & ~x[31] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[55] & ~x[56] & ~x[57] & ~x[60] & ~x[63];
			partial_clause[100] 	= partial_clause_prev[100] & ~x[9] & ~x[20] & ~x[26] & ~x[36] & ~x[39] & ~x[42];
			partial_clause[101] 	= partial_clause_prev[101] & ~x[52];
			partial_clause[102] 	= partial_clause_prev[102] & ~x[27] & ~x[58];
			partial_clause[103] 	= partial_clause_prev[103] & ~x[2] & ~x[4] & ~x[22] & ~x[24] & ~x[26] & ~x[27] & ~x[29] & ~x[32] & ~x[35] & ~x[37] & ~x[38] & ~x[49] & ~x[50] & ~x[51] & ~x[52] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[59] & ~x[60] & ~x[61];
			partial_clause[104] 	= partial_clause_prev[104] & ~x[3] & ~x[18] & ~x[23] & ~x[24] & ~x[25] & ~x[26] & ~x[29] & ~x[48] & ~x[51] & ~x[52];
			partial_clause[105] 	= partial_clause_prev[105] & ~x[0] & ~x[1] & ~x[2] & ~x[7] & ~x[9] & ~x[11] & ~x[12] & ~x[13] & ~x[27] & ~x[30] & ~x[40] & ~x[56] & ~x[63];
			partial_clause[106] 	= partial_clause_prev[106] & ~x[39];
			partial_clause[107] 	= partial_clause_prev[107] & ~x[9] & ~x[27] & ~x[28] & ~x[29] & ~x[31] & ~x[38] & ~x[39];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[2] & ~x[4] & ~x[8] & ~x[15] & ~x[33] & ~x[41] & ~x[53] & ~x[54] & ~x[56] & ~x[59] & ~x[63];
			partial_clause[109] 	= partial_clause_prev[109] & 1'b1;
			partial_clause[110] 	= partial_clause_prev[110] & ~x[41];
			partial_clause[111] 	= partial_clause_prev[111] & 1'b1;
			partial_clause[112] 	= partial_clause_prev[112] & ~x[52] & ~x[56] & ~x[63];
			partial_clause[113] 	= partial_clause_prev[113] & ~x[23] & ~x[61];
			partial_clause[114] 	= partial_clause_prev[114] & 1'b1;
			partial_clause[115] 	= partial_clause_prev[115] & ~x[0] & ~x[7] & ~x[9] & ~x[12] & ~x[33] & ~x[34] & ~x[35] & ~x[50] & ~x[55] & ~x[59] & ~x[62] & ~x[63];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[3] & ~x[6] & ~x[25] & ~x[38] & ~x[52] & ~x[59] & ~x[61];
			partial_clause[117] 	= partial_clause_prev[117] & 1'b1;
			partial_clause[118] 	= partial_clause_prev[118] & ~x[3] & ~x[8] & ~x[28] & ~x[31] & ~x[35] & ~x[57];
			partial_clause[119] 	= partial_clause_prev[119] & ~x[1] & ~x[4] & ~x[5] & ~x[29] & ~x[30] & ~x[31] & ~x[33] & ~x[35] & ~x[37] & ~x[59] & ~x[60] & ~x[62];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[1] & ~x[2] & ~x[3] & ~x[5] & ~x[6] & x[18] & ~x[27] & ~x[34] & ~x[52] & ~x[54] & ~x[55] & ~x[58] & ~x[60];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[0] & ~x[2] & ~x[24] & ~x[25] & ~x[57] & ~x[58] & ~x[61];
			partial_clause[122] 	= partial_clause_prev[122] & ~x[29] & ~x[35] & ~x[56];
			partial_clause[123] 	= partial_clause_prev[123] & ~x[4] & ~x[8] & ~x[23] & ~x[31] & ~x[33] & ~x[35] & ~x[37] & ~x[54] & ~x[57] & ~x[58] & ~x[59] & ~x[60];
			partial_clause[124] 	= partial_clause_prev[124] & ~x[25];
			partial_clause[125] 	= partial_clause_prev[125] & ~x[33] & ~x[40] & ~x[50] & ~x[54] & ~x[60];
			partial_clause[126] 	= partial_clause_prev[126] & ~x[57];
			partial_clause[127] 	= partial_clause_prev[127] & ~x[2] & ~x[4] & ~x[6] & ~x[8] & ~x[9] & ~x[27] & ~x[28] & ~x[29] & ~x[30] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[38] & ~x[59] & ~x[63];
			partial_clause[128] 	= partial_clause_prev[128] & ~x[62] & ~x[63];
			partial_clause[129] 	= partial_clause_prev[129] & ~x[8] & ~x[22] & ~x[23] & ~x[26] & ~x[28] & ~x[33] & ~x[35] & ~x[49] & ~x[51] & ~x[52] & ~x[59] & ~x[61];
			partial_clause[130] 	= partial_clause_prev[130] & ~x[3] & ~x[5] & ~x[8] & ~x[19] & ~x[51] & ~x[62];
			partial_clause[131] 	= partial_clause_prev[131] & 1'b1;
			partial_clause[132] 	= partial_clause_prev[132] & ~x[22] & ~x[28];
			partial_clause[133] 	= partial_clause_prev[133] & ~x[0] & ~x[4] & ~x[51] & ~x[52] & ~x[61];
			partial_clause[134] 	= partial_clause_prev[134] & ~x[2] & ~x[4] & ~x[6] & ~x[7] & ~x[29] & ~x[31] & ~x[33] & ~x[34] & ~x[52] & ~x[55] & ~x[62];
			partial_clause[135] 	= partial_clause_prev[135] & ~x[2] & ~x[8] & ~x[20] & ~x[29] & ~x[30] & ~x[32] & ~x[37] & ~x[52] & ~x[55];
			partial_clause[136] 	= partial_clause_prev[136] & ~x[1] & ~x[26] & ~x[28] & ~x[30] & ~x[57];
			partial_clause[137] 	= partial_clause_prev[137] & ~x[2];
			partial_clause[138] 	= partial_clause_prev[138] & 1'b1;
			partial_clause[139] 	= partial_clause_prev[139] & ~x[1] & ~x[6] & ~x[7] & ~x[35] & ~x[37] & ~x[38] & ~x[54] & ~x[58] & ~x[59] & ~x[61];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[0] & ~x[4] & ~x[24] & ~x[33] & ~x[49] & ~x[50] & ~x[51] & ~x[59] & ~x[62] & ~x[63];
			partial_clause[141] 	= partial_clause_prev[141] & ~x[6] & ~x[60];
			partial_clause[142] 	= partial_clause_prev[142] & ~x[5] & ~x[11] & ~x[32] & ~x[34] & ~x[39] & ~x[56];
			partial_clause[143] 	= partial_clause_prev[143] & ~x[2] & ~x[63];
			partial_clause[144] 	= partial_clause_prev[144] & ~x[7] & ~x[25] & ~x[32] & ~x[57] & ~x[60] & ~x[62];
			partial_clause[145] 	= partial_clause_prev[145] & 1'b1;
			partial_clause[146] 	= partial_clause_prev[146] & ~x[4] & ~x[22] & ~x[24] & ~x[52] & ~x[54] & ~x[58] & ~x[62];
			partial_clause[147] 	= partial_clause_prev[147] & ~x[4] & ~x[23] & ~x[26] & ~x[33] & ~x[34] & ~x[35] & ~x[36] & ~x[42] & ~x[55] & ~x[57];
			partial_clause[148] 	= partial_clause_prev[148] & ~x[6] & ~x[13] & ~x[31] & ~x[33] & ~x[41] & ~x[53] & ~x[59] & ~x[61] & ~x[63];
			partial_clause[149] 	= partial_clause_prev[149] & ~x[6] & ~x[34];
			partial_clause[150] 	= partial_clause_prev[150] & ~x[40] & ~x[41] & ~x[46] & ~x[48];
			partial_clause[151] 	= partial_clause_prev[151] & ~x[48];
			partial_clause[152] 	= partial_clause_prev[152] & ~x[8] & ~x[35] & ~x[54] & ~x[58];
			partial_clause[153] 	= partial_clause_prev[153] & ~x[3] & ~x[6] & ~x[36] & ~x[62];
			partial_clause[154] 	= partial_clause_prev[154] & ~x[3] & ~x[4] & ~x[24] & ~x[55] & ~x[59];
			partial_clause[155] 	= partial_clause_prev[155] & 1'b1;
			partial_clause[156] 	= partial_clause_prev[156] & 1'b1;
			partial_clause[157] 	= partial_clause_prev[157] & 1'b1;
			partial_clause[158] 	= partial_clause_prev[158] & ~x[0] & ~x[2] & ~x[4] & ~x[6] & ~x[8] & ~x[24] & ~x[25] & ~x[29] & ~x[31] & ~x[33] & ~x[34] & ~x[51] & ~x[55] & ~x[60] & ~x[63];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[27] & ~x[35] & ~x[42] & ~x[46] & ~x[50] & ~x[52] & ~x[56];
			partial_clause[160] 	= partial_clause_prev[160] & ~x[34] & ~x[38];
			partial_clause[161] 	= partial_clause_prev[161] & ~x[0] & ~x[2] & ~x[23] & ~x[26] & ~x[33] & ~x[51] & ~x[57] & ~x[62];
			partial_clause[162] 	= partial_clause_prev[162] & ~x[24] & ~x[27] & ~x[28] & ~x[31];
			partial_clause[163] 	= partial_clause_prev[163] & 1'b1;
			partial_clause[164] 	= partial_clause_prev[164] & ~x[38];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[28] & ~x[31] & ~x[63];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[7] & ~x[36] & ~x[52] & ~x[58];
			partial_clause[167] 	= partial_clause_prev[167] & ~x[47];
			partial_clause[168] 	= partial_clause_prev[168] & x[45];
			partial_clause[169] 	= partial_clause_prev[169] & 1'b1;
			partial_clause[170] 	= partial_clause_prev[170] & ~x[39];
			partial_clause[171] 	= partial_clause_prev[171] & ~x[3] & ~x[27] & ~x[57];
			partial_clause[172] 	= partial_clause_prev[172] & 1'b1;
			partial_clause[173] 	= partial_clause_prev[173] & ~x[24] & ~x[53] & ~x[57] & ~x[63];
			partial_clause[174] 	= partial_clause_prev[174] & ~x[21] & ~x[25] & ~x[26] & ~x[49] & ~x[51];
			partial_clause[175] 	= partial_clause_prev[175] & 1'b1;
			partial_clause[176] 	= partial_clause_prev[176] & ~x[20] & ~x[24];
			partial_clause[177] 	= partial_clause_prev[177] & ~x[3] & ~x[28] & ~x[50] & ~x[53] & ~x[60] & ~x[63];
			partial_clause[178] 	= partial_clause_prev[178] & ~x[38] & ~x[62];
			partial_clause[179] 	= partial_clause_prev[179] & 1'b1;
			partial_clause[180] 	= partial_clause_prev[180] & ~x[5] & x[17] & ~x[30] & ~x[54];
			partial_clause[181] 	= partial_clause_prev[181] & 1'b1;
			partial_clause[182] 	= partial_clause_prev[182] & ~x[55];
			partial_clause[183] 	= partial_clause_prev[183] & ~x[2] & ~x[5] & ~x[22] & ~x[24] & ~x[25] & ~x[26] & ~x[28] & ~x[29] & ~x[31] & ~x[33] & ~x[51] & ~x[52] & ~x[55] & ~x[59] & ~x[60] & ~x[63];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[6] & ~x[8] & ~x[22] & ~x[26] & ~x[35] & ~x[58];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[1] & ~x[11] & ~x[13] & ~x[15] & ~x[16] & ~x[17] & ~x[43] & ~x[50];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[36] & ~x[38] & ~x[40] & ~x[54] & ~x[55] & ~x[57];
			partial_clause[187] 	= partial_clause_prev[187] & ~x[1] & ~x[5] & ~x[6] & ~x[12] & ~x[30] & ~x[31] & ~x[34] & ~x[38] & ~x[58];
			partial_clause[188] 	= partial_clause_prev[188] & ~x[7] & ~x[60];
			partial_clause[189] 	= partial_clause_prev[189] & 1'b1;
			partial_clause[190] 	= partial_clause_prev[190] & ~x[3] & ~x[5] & ~x[8] & ~x[31] & ~x[33] & ~x[55] & ~x[59];
			partial_clause[191] 	= partial_clause_prev[191] & ~x[2] & ~x[20] & ~x[33] & ~x[38] & ~x[54] & ~x[63];
			partial_clause[192] 	= partial_clause_prev[192] & ~x[1] & ~x[2] & ~x[40];
			partial_clause[193] 	= partial_clause_prev[193] & ~x[0] & ~x[4] & ~x[10] & ~x[12] & ~x[27] & ~x[37] & ~x[55];
			partial_clause[194] 	= partial_clause_prev[194] & ~x[3] & ~x[5] & ~x[7];
			partial_clause[195] 	= partial_clause_prev[195] & ~x[0] & ~x[3] & ~x[5] & ~x[6] & ~x[20] & ~x[21] & ~x[22] & ~x[31] & ~x[33] & ~x[48] & ~x[49] & ~x[54] & ~x[61];
			partial_clause[196] 	= partial_clause_prev[196] & 1'b1;
			partial_clause[197] 	= partial_clause_prev[197] & ~x[0] & ~x[5] & ~x[6] & ~x[7] & ~x[37] & ~x[41] & ~x[44] & ~x[53] & ~x[56] & ~x[57] & ~x[58] & ~x[61];
			partial_clause[198] 	= partial_clause_prev[198] & 1'b1;
			partial_clause[199] 	= partial_clause_prev[199] & ~x[49] & ~x[52];
			partial_clause[200] 	= partial_clause_prev[200] & ~x[5] & ~x[54] & ~x[60] & ~x[61];
			partial_clause[201] 	= partial_clause_prev[201] & ~x[5] & ~x[20] & ~x[24] & ~x[25] & ~x[59] & ~x[63];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[4] & ~x[5] & ~x[8] & ~x[9] & ~x[26] & ~x[38] & ~x[39] & ~x[44] & ~x[51] & ~x[53] & ~x[63];
			partial_clause[203] 	= partial_clause_prev[203] & ~x[23] & ~x[32];
			partial_clause[204] 	= partial_clause_prev[204] & ~x[13] & ~x[28] & ~x[31] & ~x[36] & ~x[41] & ~x[42] & ~x[58] & ~x[59];
			partial_clause[205] 	= partial_clause_prev[205] & ~x[51];
			partial_clause[206] 	= partial_clause_prev[206] & ~x[0] & ~x[1] & ~x[2] & x[16] & ~x[27] & ~x[29] & ~x[31] & ~x[34] & ~x[37] & ~x[52] & ~x[63];
			partial_clause[207] 	= partial_clause_prev[207] & ~x[11] & ~x[39] & ~x[41] & ~x[51];
			partial_clause[208] 	= partial_clause_prev[208] & ~x[0] & ~x[35] & ~x[56] & ~x[57];
			partial_clause[209] 	= partial_clause_prev[209] & 1'b1;
			partial_clause[210] 	= partial_clause_prev[210] & ~x[0] & ~x[2] & ~x[25] & ~x[27] & ~x[29] & ~x[32] & ~x[33] & ~x[34] & ~x[48];
			partial_clause[211] 	= partial_clause_prev[211] & 1'b1;
			partial_clause[212] 	= partial_clause_prev[212] & ~x[32] & ~x[38] & ~x[44] & ~x[50];
			partial_clause[213] 	= partial_clause_prev[213] & 1'b1;
			partial_clause[214] 	= partial_clause_prev[214] & ~x[3] & ~x[15] & ~x[21] & ~x[46];
			partial_clause[215] 	= partial_clause_prev[215] & ~x[48] & ~x[49];
			partial_clause[216] 	= partial_clause_prev[216] & ~x[5];
			partial_clause[217] 	= partial_clause_prev[217] & ~x[0] & ~x[9] & ~x[10] & ~x[29] & ~x[32] & ~x[41] & ~x[49];
			partial_clause[218] 	= partial_clause_prev[218] & 1'b1;
			partial_clause[219] 	= partial_clause_prev[219] & ~x[13] & ~x[15] & ~x[18] & ~x[19] & ~x[20] & ~x[22] & ~x[44];
			partial_clause[220] 	= partial_clause_prev[220] & ~x[0] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[24] & ~x[31] & ~x[33] & ~x[36] & ~x[38] & ~x[51] & ~x[52] & ~x[56] & ~x[58] & ~x[61];
			partial_clause[221] 	= partial_clause_prev[221] & 1'b1;
			partial_clause[222] 	= partial_clause_prev[222] & 1'b1;
			partial_clause[223] 	= partial_clause_prev[223] & ~x[3];
			partial_clause[224] 	= partial_clause_prev[224] & ~x[5] & ~x[6] & ~x[28] & ~x[34] & ~x[35] & ~x[37] & ~x[40] & ~x[41] & ~x[50] & ~x[54] & ~x[56] & ~x[57];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[54] & ~x[56] & ~x[60];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[0] & ~x[1] & ~x[3] & ~x[7] & ~x[12] & ~x[15] & ~x[27] & ~x[28] & ~x[36] & ~x[38] & ~x[40] & ~x[42] & ~x[58] & ~x[59] & ~x[61];
			partial_clause[227] 	= partial_clause_prev[227] & ~x[1] & ~x[6] & ~x[17] & ~x[29] & ~x[33] & ~x[41] & ~x[42] & ~x[44] & ~x[59] & ~x[63];
			partial_clause[228] 	= partial_clause_prev[228] & ~x[0] & ~x[6] & ~x[29] & ~x[54] & ~x[57] & ~x[58] & ~x[59];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[0] & ~x[9] & ~x[25] & ~x[27] & ~x[33] & ~x[36] & ~x[40] & ~x[52] & ~x[53] & ~x[59];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[3] & ~x[5] & ~x[6] & ~x[7] & ~x[27] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[37] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[231] 	= partial_clause_prev[231] & ~x[1] & ~x[27] & ~x[42] & ~x[58];
			partial_clause[232] 	= partial_clause_prev[232] & 1'b1;
			partial_clause[233] 	= partial_clause_prev[233] & 1'b1;
			partial_clause[234] 	= partial_clause_prev[234] & ~x[3] & ~x[17] & ~x[20] & ~x[38];
			partial_clause[235] 	= partial_clause_prev[235] & 1'b1;
			partial_clause[236] 	= partial_clause_prev[236] & ~x[30];
			partial_clause[237] 	= partial_clause_prev[237] & ~x[28] & ~x[58];
			partial_clause[238] 	= partial_clause_prev[238] & 1'b1;
			partial_clause[239] 	= partial_clause_prev[239] & ~x[5] & ~x[51];
			partial_clause[240] 	= partial_clause_prev[240] & ~x[0] & ~x[25] & ~x[28] & ~x[35] & ~x[51] & ~x[62];
			partial_clause[241] 	= partial_clause_prev[241] & ~x[7] & ~x[59];
			partial_clause[242] 	= partial_clause_prev[242] & ~x[5] & ~x[6] & ~x[24] & ~x[25] & ~x[30] & ~x[55] & ~x[56] & ~x[57] & ~x[59];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[2] & ~x[10] & ~x[26] & ~x[27] & ~x[39] & ~x[56] & ~x[61];
			partial_clause[244] 	= partial_clause_prev[244] & ~x[6];
			partial_clause[245] 	= partial_clause_prev[245] & 1'b1;
			partial_clause[246] 	= partial_clause_prev[246] & 1'b1;
			partial_clause[247] 	= partial_clause_prev[247] & ~x[2] & ~x[3] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[25] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[38] & ~x[51] & ~x[63];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[0] & ~x[4] & ~x[6] & ~x[10] & ~x[11] & ~x[13] & ~x[25] & ~x[29] & ~x[32] & ~x[34] & ~x[35] & ~x[38] & ~x[45] & ~x[58] & ~x[60] & ~x[63];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[0];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[1] & ~x[6] & ~x[10] & ~x[25] & ~x[26] & ~x[28] & ~x[31] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[38] & ~x[51] & ~x[54] & ~x[56] & ~x[57] & ~x[58];
			partial_clause[251] 	= partial_clause_prev[251] & 1'b1;
			partial_clause[252] 	= partial_clause_prev[252] & ~x[0] & ~x[2] & ~x[4] & ~x[7] & ~x[11] & ~x[12] & ~x[36] & ~x[37] & ~x[54] & ~x[57] & ~x[61];
			partial_clause[253] 	= partial_clause_prev[253] & ~x[35];
			partial_clause[254] 	= partial_clause_prev[254] & ~x[4] & ~x[5] & ~x[23] & ~x[33] & ~x[34] & ~x[52];
			partial_clause[255] 	= partial_clause_prev[255] & ~x[16] & ~x[19] & ~x[23] & ~x[25] & ~x[26] & ~x[39] & ~x[46] & ~x[47] & ~x[49];
			partial_clause[256] 	= partial_clause_prev[256] & 1'b1;
			partial_clause[257] 	= partial_clause_prev[257] & ~x[25] & ~x[33];
			partial_clause[258] 	= partial_clause_prev[258] & ~x[5] & ~x[29] & ~x[30] & ~x[31] & ~x[60];
			partial_clause[259] 	= partial_clause_prev[259] & 1'b1;
			partial_clause[260] 	= partial_clause_prev[260] & ~x[3] & ~x[6] & ~x[10] & ~x[28] & ~x[57];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[1] & ~x[6] & ~x[23] & ~x[34] & ~x[58];
			partial_clause[262] 	= partial_clause_prev[262] & ~x[30];
			partial_clause[263] 	= partial_clause_prev[263] & ~x[5] & ~x[24] & ~x[50];
			partial_clause[264] 	= partial_clause_prev[264] & ~x[0] & ~x[3] & ~x[35];
			partial_clause[265] 	= partial_clause_prev[265] & 1'b1;
			partial_clause[266] 	= partial_clause_prev[266] & ~x[1] & ~x[22] & ~x[25] & ~x[31] & ~x[34] & ~x[37] & ~x[41] & ~x[54] & ~x[60];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[2] & ~x[6] & ~x[22] & ~x[25] & ~x[26] & ~x[27] & ~x[34] & ~x[35] & ~x[52] & ~x[53] & ~x[54] & ~x[59] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[1] & ~x[5] & ~x[7] & ~x[10] & ~x[28] & ~x[29] & ~x[33] & ~x[40] & ~x[58] & ~x[59] & ~x[60] & ~x[62];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[4] & ~x[5] & ~x[6] & ~x[21] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[27] & ~x[29] & ~x[30] & ~x[35] & ~x[36] & ~x[38] & ~x[39] & ~x[40] & ~x[41] & ~x[42] & ~x[46] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[52] & ~x[54] & ~x[55] & ~x[57] & ~x[58] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[270] 	= partial_clause_prev[270] & 1'b1;
			partial_clause[271] 	= partial_clause_prev[271] & ~x[0] & ~x[7] & ~x[33] & ~x[55];
			partial_clause[272] 	= partial_clause_prev[272] & ~x[1] & ~x[3] & ~x[31] & ~x[32] & ~x[58];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[0] & ~x[1] & ~x[2] & ~x[6] & ~x[7] & ~x[8] & ~x[11] & ~x[12] & ~x[14] & ~x[15] & ~x[29] & ~x[30] & ~x[32] & ~x[35] & ~x[40] & ~x[42] & ~x[47] & ~x[60] & ~x[61] & ~x[63];
			partial_clause[274] 	= partial_clause_prev[274] & ~x[7] & ~x[55] & ~x[63];
			partial_clause[275] 	= partial_clause_prev[275] & ~x[40];
			partial_clause[276] 	= partial_clause_prev[276] & ~x[6] & ~x[48];
			partial_clause[277] 	= partial_clause_prev[277] & ~x[24] & ~x[25] & ~x[28] & ~x[56] & ~x[57] & ~x[63];
			partial_clause[278] 	= partial_clause_prev[278] & 1'b1;
			partial_clause[279] 	= partial_clause_prev[279] & ~x[4] & ~x[8] & ~x[13] & ~x[33] & ~x[35] & ~x[41] & ~x[42];
			partial_clause[280] 	= partial_clause_prev[280] & 1'b1;
			partial_clause[281] 	= partial_clause_prev[281] & ~x[7] & ~x[8] & ~x[11] & ~x[42] & ~x[49] & ~x[58] & ~x[60] & ~x[63];
			partial_clause[282] 	= partial_clause_prev[282] & ~x[28] & ~x[31] & ~x[34] & ~x[55] & ~x[57];
			partial_clause[283] 	= partial_clause_prev[283] & ~x[4] & ~x[11] & ~x[18] & ~x[47];
			partial_clause[284] 	= partial_clause_prev[284] & 1'b1;
			partial_clause[285] 	= partial_clause_prev[285] & 1'b1;
			partial_clause[286] 	= partial_clause_prev[286] & ~x[20] & ~x[21];
			partial_clause[287] 	= partial_clause_prev[287] & ~x[0] & ~x[2] & ~x[6] & ~x[10] & ~x[23] & ~x[28] & ~x[29] & ~x[30] & ~x[31] & ~x[32] & ~x[36] & ~x[38] & ~x[49] & ~x[51] & ~x[58] & ~x[59];
			partial_clause[288] 	= partial_clause_prev[288] & ~x[9] & ~x[51];
			partial_clause[289] 	= partial_clause_prev[289] & ~x[1] & ~x[7] & ~x[32] & ~x[63];
			partial_clause[290] 	= partial_clause_prev[290] & ~x[3] & ~x[4] & ~x[8] & ~x[13] & ~x[33] & ~x[37];
			partial_clause[291] 	= partial_clause_prev[291] & 1'b1;
			partial_clause[292] 	= partial_clause_prev[292] & ~x[1] & ~x[3] & ~x[36] & ~x[48] & ~x[49] & ~x[59];
			partial_clause[293] 	= partial_clause_prev[293] & ~x[7] & ~x[34] & ~x[63];
			partial_clause[294] 	= partial_clause_prev[294] & ~x[2] & ~x[10] & ~x[11] & ~x[12] & ~x[17];
			partial_clause[295] 	= partial_clause_prev[295] & ~x[29] & ~x[37];
			partial_clause[296] 	= partial_clause_prev[296] & 1'b1;
			partial_clause[297] 	= partial_clause_prev[297] & ~x[5] & ~x[48] & ~x[51];
			partial_clause[298] 	= partial_clause_prev[298] & 1'b1;
			partial_clause[299] 	= partial_clause_prev[299] & ~x[6] & ~x[36] & ~x[54] & ~x[55] & ~x[56];
			partial_clause[300] 	= partial_clause_prev[300] & ~x[23] & ~x[36] & ~x[53] & ~x[60];
			partial_clause[301] 	= partial_clause_prev[301] & ~x[7] & ~x[24] & ~x[48] & ~x[51] & ~x[54] & ~x[55];
			partial_clause[302] 	= partial_clause_prev[302] & ~x[7] & ~x[31];
			partial_clause[303] 	= partial_clause_prev[303] & ~x[3] & ~x[52] & ~x[63];
			partial_clause[304] 	= partial_clause_prev[304] & ~x[51];
			partial_clause[305] 	= partial_clause_prev[305] & ~x[26] & ~x[63];
			partial_clause[306] 	= partial_clause_prev[306] & ~x[55];
			partial_clause[307] 	= partial_clause_prev[307] & ~x[3] & ~x[8] & ~x[32] & ~x[35] & ~x[36] & ~x[47];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[0] & ~x[8] & ~x[9] & ~x[11] & ~x[26] & ~x[29] & ~x[31] & ~x[39];
			partial_clause[309] 	= partial_clause_prev[309] & ~x[2] & ~x[32] & ~x[35] & ~x[37] & ~x[53] & ~x[57] & ~x[63];
			partial_clause[310] 	= partial_clause_prev[310] & 1'b1;
			partial_clause[311] 	= partial_clause_prev[311] & ~x[9] & ~x[22] & ~x[47] & ~x[50] & ~x[51];
			partial_clause[312] 	= partial_clause_prev[312] & ~x[5];
			partial_clause[313] 	= partial_clause_prev[313] & ~x[14];
			partial_clause[314] 	= partial_clause_prev[314] & ~x[28] & ~x[37] & ~x[55];
			partial_clause[315] 	= partial_clause_prev[315] & ~x[2] & ~x[5] & ~x[9] & ~x[10] & ~x[30] & ~x[33] & ~x[51] & ~x[61] & ~x[63];
			partial_clause[316] 	= partial_clause_prev[316] & ~x[1] & ~x[3] & ~x[5] & ~x[27] & ~x[28] & ~x[29] & ~x[34] & ~x[36] & ~x[59];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[6] & ~x[32] & ~x[36] & ~x[38] & ~x[47] & ~x[59] & ~x[63];
			partial_clause[318] 	= partial_clause_prev[318] & ~x[21] & ~x[25] & ~x[35] & ~x[61];
			partial_clause[319] 	= partial_clause_prev[319] & ~x[32];
			partial_clause[320] 	= partial_clause_prev[320] & ~x[5] & ~x[12] & ~x[13] & ~x[14] & ~x[26] & ~x[29] & ~x[35] & ~x[36] & ~x[37] & ~x[44] & ~x[45] & ~x[47] & ~x[48] & ~x[56];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[8] & ~x[31] & ~x[54] & ~x[59] & ~x[60];
			partial_clause[322] 	= partial_clause_prev[322] & ~x[48] & ~x[50] & ~x[58];
			partial_clause[323] 	= partial_clause_prev[323] & ~x[9] & ~x[59];
			partial_clause[324] 	= partial_clause_prev[324] & ~x[4] & ~x[36];
			partial_clause[325] 	= partial_clause_prev[325] & ~x[1] & ~x[3] & ~x[7] & ~x[21] & ~x[23] & ~x[25] & ~x[29] & ~x[34] & ~x[35] & ~x[37] & ~x[42] & ~x[48] & ~x[49] & ~x[50] & ~x[52] & ~x[53] & ~x[54] & ~x[57] & ~x[58] & ~x[63];
			partial_clause[326] 	= partial_clause_prev[326] & ~x[2] & ~x[5] & ~x[9] & ~x[10] & ~x[27] & ~x[30] & ~x[35] & ~x[36] & ~x[56];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[1] & ~x[6] & ~x[11] & ~x[13] & ~x[22] & ~x[25] & ~x[27] & ~x[33] & ~x[55];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[5] & ~x[9] & ~x[22] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[41];
			partial_clause[329] 	= partial_clause_prev[329] & ~x[51];
			partial_clause[330] 	= partial_clause_prev[330] & ~x[1] & ~x[6] & ~x[34] & ~x[37] & ~x[61];
			partial_clause[331] 	= partial_clause_prev[331] & ~x[0] & ~x[4] & ~x[23] & ~x[31] & ~x[50] & ~x[54] & ~x[58];
			partial_clause[332] 	= partial_clause_prev[332] & ~x[8] & ~x[32] & ~x[57];
			partial_clause[333] 	= partial_clause_prev[333] & ~x[2] & ~x[36];
			partial_clause[334] 	= partial_clause_prev[334] & ~x[0];
			partial_clause[335] 	= partial_clause_prev[335] & 1'b1;
			partial_clause[336] 	= partial_clause_prev[336] & ~x[25];
			partial_clause[337] 	= partial_clause_prev[337] & ~x[3] & ~x[5] & ~x[9] & ~x[17] & ~x[20] & ~x[37] & ~x[39] & ~x[43] & ~x[44] & ~x[45] & ~x[50] & ~x[58];
			partial_clause[338] 	= partial_clause_prev[338] & ~x[14] & ~x[19];
			partial_clause[339] 	= partial_clause_prev[339] & ~x[5] & ~x[26] & ~x[28] & ~x[31] & ~x[35] & ~x[50] & ~x[56];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[2] & ~x[28] & ~x[31] & ~x[32] & ~x[36] & ~x[55] & ~x[58] & ~x[61] & ~x[62];
			partial_clause[341] 	= partial_clause_prev[341] & 1'b1;
			partial_clause[342] 	= partial_clause_prev[342] & ~x[4] & ~x[5] & ~x[28] & ~x[32] & ~x[33] & ~x[60];
			partial_clause[343] 	= partial_clause_prev[343] & ~x[1] & ~x[4] & ~x[22] & ~x[27] & ~x[35] & ~x[36] & ~x[49] & ~x[53] & ~x[55] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[8];
			partial_clause[345] 	= partial_clause_prev[345] & ~x[31] & ~x[33] & ~x[54];
			partial_clause[346] 	= partial_clause_prev[346] & 1'b1;
			partial_clause[347] 	= partial_clause_prev[347] & ~x[3] & ~x[28] & ~x[50] & ~x[60];
			partial_clause[348] 	= partial_clause_prev[348] & ~x[1] & ~x[5] & ~x[40];
			partial_clause[349] 	= partial_clause_prev[349] & ~x[33];
			partial_clause[350] 	= partial_clause_prev[350] & ~x[1] & ~x[3] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[12] & ~x[27] & ~x[28] & ~x[32] & ~x[33] & ~x[38] & ~x[42] & ~x[54] & ~x[56] & ~x[57] & ~x[58] & ~x[60] & ~x[61];
			partial_clause[351] 	= partial_clause_prev[351] & ~x[38] & ~x[59];
			partial_clause[352] 	= partial_clause_prev[352] & 1'b1;
			partial_clause[353] 	= partial_clause_prev[353] & 1'b1;
			partial_clause[354] 	= partial_clause_prev[354] & ~x[40] & ~x[41] & ~x[47] & ~x[53] & ~x[56] & ~x[62];
			partial_clause[355] 	= partial_clause_prev[355] & ~x[32] & ~x[34] & ~x[38] & ~x[40];
			partial_clause[356] 	= partial_clause_prev[356] & ~x[27] & ~x[53] & ~x[59] & ~x[63];
			partial_clause[357] 	= partial_clause_prev[357] & 1'b1;
			partial_clause[358] 	= partial_clause_prev[358] & ~x[5] & ~x[9] & ~x[31] & ~x[34] & ~x[37] & ~x[39] & ~x[57];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[27] & ~x[35] & ~x[58];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[4] & ~x[8] & ~x[9] & ~x[29] & ~x[31] & ~x[37] & ~x[39] & ~x[57] & ~x[59] & ~x[61];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[7] & ~x[8];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[10] & ~x[21] & ~x[33] & ~x[50];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[7] & ~x[8] & ~x[11] & ~x[12] & ~x[23] & ~x[26] & ~x[32] & ~x[33] & ~x[39] & ~x[52] & ~x[53] & ~x[59] & ~x[60];
			partial_clause[364] 	= partial_clause_prev[364] & ~x[17] & ~x[18] & ~x[19] & ~x[37] & ~x[41] & ~x[42] & ~x[45] & ~x[58] & ~x[60];
			partial_clause[365] 	= partial_clause_prev[365] & ~x[58];
			partial_clause[366] 	= partial_clause_prev[366] & ~x[28] & ~x[29] & ~x[33] & ~x[35] & ~x[55] & ~x[61];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[0] & ~x[27] & ~x[35] & ~x[36] & ~x[45] & ~x[51];
			partial_clause[368] 	= partial_clause_prev[368] & 1'b1;
			partial_clause[369] 	= partial_clause_prev[369] & ~x[2] & ~x[8] & ~x[10] & ~x[31];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[9] & ~x[10] & ~x[12] & ~x[23] & ~x[24] & ~x[25] & ~x[54] & ~x[58];
			partial_clause[371] 	= partial_clause_prev[371] & ~x[10] & ~x[25] & ~x[39] & ~x[45];
			partial_clause[372] 	= partial_clause_prev[372] & ~x[25] & ~x[31];
			partial_clause[373] 	= partial_clause_prev[373] & 1'b1;
			partial_clause[374] 	= partial_clause_prev[374] & 1'b1;
			partial_clause[375] 	= partial_clause_prev[375] & ~x[50];
			partial_clause[376] 	= partial_clause_prev[376] & ~x[0] & ~x[2] & ~x[8] & ~x[9] & ~x[12] & ~x[14] & ~x[34] & ~x[56] & ~x[58];
			partial_clause[377] 	= partial_clause_prev[377] & 1'b1;
			partial_clause[378] 	= partial_clause_prev[378] & ~x[5] & ~x[31] & ~x[34] & ~x[36] & ~x[62];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[27] & ~x[58];
			partial_clause[380] 	= partial_clause_prev[380] & 1'b1;
			partial_clause[381] 	= partial_clause_prev[381] & ~x[1] & ~x[11] & ~x[12] & ~x[32] & ~x[37] & ~x[42] & ~x[43] & ~x[44] & ~x[45] & ~x[47] & ~x[48] & ~x[51] & ~x[53] & ~x[55] & ~x[59] & ~x[62];
			partial_clause[382] 	= partial_clause_prev[382] & 1'b1;
			partial_clause[383] 	= partial_clause_prev[383] & 1'b1;
			partial_clause[384] 	= partial_clause_prev[384] & 1'b1;
			partial_clause[385] 	= partial_clause_prev[385] & ~x[58];
			partial_clause[386] 	= partial_clause_prev[386] & ~x[6] & ~x[42];
			partial_clause[387] 	= partial_clause_prev[387] & ~x[8] & ~x[9] & ~x[10] & ~x[28] & ~x[33] & ~x[56] & ~x[58] & ~x[59] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[1] & ~x[4] & ~x[7] & ~x[29] & ~x[33] & ~x[34] & ~x[37] & ~x[39] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[60] & ~x[61];
			partial_clause[389] 	= partial_clause_prev[389] & 1'b1;
			partial_clause[390] 	= partial_clause_prev[390] & ~x[5] & ~x[8] & ~x[28] & ~x[30] & ~x[32] & ~x[34] & ~x[56] & ~x[61];
			partial_clause[391] 	= partial_clause_prev[391] & 1'b1;
			partial_clause[392] 	= partial_clause_prev[392] & ~x[20] & ~x[48];
			partial_clause[393] 	= partial_clause_prev[393] & ~x[56];
			partial_clause[394] 	= partial_clause_prev[394] & ~x[34] & ~x[55];
			partial_clause[395] 	= partial_clause_prev[395] & ~x[38];
			partial_clause[396] 	= partial_clause_prev[396] & ~x[26];
			partial_clause[397] 	= partial_clause_prev[397] & ~x[0];
			partial_clause[398] 	= partial_clause_prev[398] & 1'b1;
			partial_clause[399] 	= partial_clause_prev[399] & ~x[49];
			partial_clause[400] 	= partial_clause_prev[400] & ~x[1] & ~x[3] & ~x[7] & ~x[8] & ~x[9] & ~x[10] & ~x[38];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[3] & ~x[9] & ~x[20] & ~x[21] & ~x[25] & ~x[32] & ~x[37] & ~x[53] & ~x[55] & ~x[56];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[0] & ~x[26] & ~x[38] & ~x[51] & ~x[52] & ~x[59];
			partial_clause[403] 	= partial_clause_prev[403] & ~x[12] & ~x[28] & ~x[38] & ~x[61] & ~x[62];
			partial_clause[404] 	= partial_clause_prev[404] & 1'b1;
			partial_clause[405] 	= partial_clause_prev[405] & ~x[0] & ~x[3] & ~x[24] & ~x[52];
			partial_clause[406] 	= partial_clause_prev[406] & ~x[33] & ~x[47] & ~x[55];
			partial_clause[407] 	= partial_clause_prev[407] & ~x[60];
			partial_clause[408] 	= partial_clause_prev[408] & ~x[24];
			partial_clause[409] 	= partial_clause_prev[409] & ~x[0] & ~x[2] & ~x[3] & ~x[4] & ~x[6] & ~x[10] & ~x[11] & ~x[21] & ~x[23] & ~x[24] & ~x[26] & ~x[32] & ~x[33] & ~x[39] & ~x[41] & ~x[42] & ~x[49] & ~x[50] & ~x[52] & ~x[53] & ~x[54] & ~x[56] & ~x[57] & ~x[59] & ~x[60] & ~x[61];
			partial_clause[410] 	= partial_clause_prev[410] & ~x[25] & ~x[28] & ~x[53] & ~x[61];
			partial_clause[411] 	= partial_clause_prev[411] & ~x[4] & ~x[14] & ~x[15] & ~x[31] & ~x[35] & ~x[43];
			partial_clause[412] 	= partial_clause_prev[412] & ~x[9] & ~x[35] & ~x[36] & ~x[50] & ~x[53] & ~x[54];
			partial_clause[413] 	= partial_clause_prev[413] & ~x[0] & ~x[10] & ~x[26] & ~x[30] & ~x[57];
			partial_clause[414] 	= partial_clause_prev[414] & ~x[22] & ~x[24] & ~x[31];
			partial_clause[415] 	= partial_clause_prev[415] & ~x[6] & ~x[29] & ~x[30] & ~x[62];
			partial_clause[416] 	= partial_clause_prev[416] & ~x[0] & ~x[1] & ~x[3] & ~x[22] & ~x[26] & ~x[37] & ~x[38] & ~x[39] & ~x[41] & ~x[48] & ~x[50] & ~x[51] & ~x[55] & ~x[57] & ~x[60] & ~x[61];
			partial_clause[417] 	= partial_clause_prev[417] & x[15] & ~x[23] & ~x[31] & ~x[51];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[8] & ~x[11] & ~x[26] & ~x[31] & ~x[41] & ~x[60] & ~x[61];
			partial_clause[419] 	= partial_clause_prev[419] & 1'b1;
			partial_clause[420] 	= partial_clause_prev[420] & 1'b1;
			partial_clause[421] 	= partial_clause_prev[421] & ~x[9] & ~x[28] & ~x[32];
			partial_clause[422] 	= partial_clause_prev[422] & ~x[5] & ~x[32] & ~x[34] & ~x[59];
			partial_clause[423] 	= partial_clause_prev[423] & ~x[37] & ~x[60];
			partial_clause[424] 	= partial_clause_prev[424] & ~x[6];
			partial_clause[425] 	= partial_clause_prev[425] & ~x[1];
			partial_clause[426] 	= partial_clause_prev[426] & ~x[3] & ~x[5] & ~x[6] & ~x[7] & x[17] & ~x[25] & ~x[29] & ~x[32] & ~x[35] & ~x[52] & ~x[54] & ~x[55] & ~x[63];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[7] & ~x[25] & ~x[27] & ~x[61] & ~x[62];
			partial_clause[428] 	= partial_clause_prev[428] & ~x[14] & ~x[23] & ~x[24] & ~x[25] & ~x[44];
			partial_clause[429] 	= partial_clause_prev[429] & 1'b1;
			partial_clause[430] 	= partial_clause_prev[430] & ~x[1] & ~x[3] & ~x[24] & ~x[26] & ~x[30] & ~x[33] & ~x[62];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[0] & ~x[31] & ~x[57] & ~x[61] & ~x[62];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[0] & ~x[25] & ~x[31] & ~x[32] & ~x[33] & ~x[34] & ~x[52] & ~x[56] & ~x[58] & ~x[59] & ~x[63];
			partial_clause[433] 	= partial_clause_prev[433] & ~x[28] & ~x[32] & ~x[54] & ~x[56];
			partial_clause[434] 	= partial_clause_prev[434] & 1'b1;
			partial_clause[435] 	= partial_clause_prev[435] & ~x[0] & ~x[2] & ~x[4] & ~x[5] & ~x[25] & ~x[26] & ~x[27] & ~x[51] & ~x[52] & ~x[54] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[2] & ~x[5] & ~x[34];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[4] & ~x[24] & ~x[27] & ~x[29] & ~x[30] & ~x[31] & ~x[35] & ~x[37] & ~x[47] & ~x[49] & ~x[50] & ~x[51] & ~x[53] & ~x[59] & ~x[62];
			partial_clause[438] 	= partial_clause_prev[438] & ~x[58];
			partial_clause[439] 	= partial_clause_prev[439] & ~x[0] & ~x[5] & ~x[8] & ~x[38];
			partial_clause[440] 	= partial_clause_prev[440] & ~x[8] & ~x[43] & ~x[58];
			partial_clause[441] 	= partial_clause_prev[441] & ~x[57];
			partial_clause[442] 	= partial_clause_prev[442] & 1'b1;
			partial_clause[443] 	= partial_clause_prev[443] & ~x[4] & ~x[23] & ~x[29] & ~x[54] & ~x[59];
			partial_clause[444] 	= partial_clause_prev[444] & 1'b1;
			partial_clause[445] 	= partial_clause_prev[445] & 1'b1;
			partial_clause[446] 	= partial_clause_prev[446] & ~x[35] & ~x[55];
			partial_clause[447] 	= partial_clause_prev[447] & x[14] & ~x[55] & ~x[61];
			partial_clause[448] 	= partial_clause_prev[448] & 1'b1;
			partial_clause[449] 	= partial_clause_prev[449] & ~x[1] & ~x[2] & ~x[34] & ~x[37] & ~x[57];
			partial_clause[450] 	= partial_clause_prev[450] & ~x[10] & ~x[46] & ~x[57] & ~x[58];
			partial_clause[451] 	= partial_clause_prev[451] & 1'b1;
			partial_clause[452] 	= partial_clause_prev[452] & 1'b1;
			partial_clause[453] 	= partial_clause_prev[453] & ~x[0] & ~x[43];
			partial_clause[454] 	= partial_clause_prev[454] & ~x[29] & ~x[34] & ~x[47] & ~x[49] & ~x[56] & ~x[59] & ~x[60] & ~x[63];
			partial_clause[455] 	= partial_clause_prev[455] & ~x[8] & ~x[9] & ~x[30] & ~x[33] & ~x[35] & ~x[36];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[0] & ~x[1] & ~x[5] & ~x[7] & ~x[8] & ~x[22] & ~x[23] & ~x[24] & ~x[28] & ~x[29] & ~x[30] & ~x[35] & ~x[37] & ~x[47];
			partial_clause[457] 	= partial_clause_prev[457] & 1'b1;
			partial_clause[458] 	= partial_clause_prev[458] & ~x[2] & ~x[23] & ~x[24] & ~x[26] & ~x[27] & ~x[28] & ~x[34] & ~x[56];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[0] & ~x[6] & ~x[9] & ~x[37] & ~x[38] & ~x[39] & ~x[48] & ~x[49] & ~x[52];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[0] & ~x[1] & ~x[7] & ~x[36] & ~x[49] & ~x[51] & ~x[61];
			partial_clause[461] 	= partial_clause_prev[461] & ~x[8] & ~x[11] & ~x[59];
			partial_clause[462] 	= partial_clause_prev[462] & ~x[2] & ~x[55];
			partial_clause[463] 	= partial_clause_prev[463] & ~x[24];
			partial_clause[464] 	= partial_clause_prev[464] & ~x[37] & ~x[52];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[5] & ~x[6] & ~x[8] & ~x[29] & ~x[34] & ~x[35] & ~x[36] & ~x[57] & ~x[63];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[2] & ~x[4] & ~x[8] & ~x[12] & ~x[26] & ~x[31] & ~x[33] & ~x[34] & ~x[40] & ~x[49] & ~x[62];
			partial_clause[467] 	= partial_clause_prev[467] & ~x[41] & ~x[62];
			partial_clause[468] 	= partial_clause_prev[468] & ~x[21] & ~x[34] & ~x[46] & ~x[49] & ~x[50] & ~x[53] & ~x[56] & ~x[58];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[9] & ~x[12] & ~x[24] & ~x[29] & ~x[32] & ~x[38];
			partial_clause[470] 	= partial_clause_prev[470] & ~x[59];
			partial_clause[471] 	= partial_clause_prev[471] & ~x[3] & ~x[5] & ~x[7] & ~x[21] & ~x[24] & ~x[27] & ~x[29] & ~x[31] & ~x[33] & ~x[38] & ~x[56];
			partial_clause[472] 	= partial_clause_prev[472] & ~x[34] & ~x[55];
			partial_clause[473] 	= partial_clause_prev[473] & ~x[1] & ~x[2] & ~x[24] & ~x[26] & ~x[35] & ~x[53] & ~x[60];
			partial_clause[474] 	= partial_clause_prev[474] & ~x[18] & ~x[33] & ~x[47];
			partial_clause[475] 	= partial_clause_prev[475] & ~x[10] & ~x[25] & ~x[60] & ~x[62];
			partial_clause[476] 	= partial_clause_prev[476] & ~x[15] & ~x[16] & ~x[28] & ~x[29] & ~x[31] & ~x[63];
			partial_clause[477] 	= partial_clause_prev[477] & ~x[5] & ~x[30] & ~x[41] & ~x[50] & ~x[51] & ~x[57] & ~x[60] & ~x[61];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[0] & ~x[6] & ~x[9] & ~x[23] & ~x[34] & ~x[35] & ~x[37] & ~x[42] & ~x[49] & ~x[52];
			partial_clause[479] 	= partial_clause_prev[479] & ~x[18] & ~x[44];
			partial_clause[480] 	= partial_clause_prev[480] & ~x[0] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[27] & ~x[29] & ~x[30] & ~x[32] & ~x[33] & ~x[34] & ~x[35] & ~x[36] & ~x[38] & ~x[52] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[59] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[481] 	= partial_clause_prev[481] & ~x[4] & ~x[38] & ~x[60];
			partial_clause[482] 	= partial_clause_prev[482] & ~x[8] & ~x[29] & ~x[35] & ~x[55] & ~x[57];
			partial_clause[483] 	= partial_clause_prev[483] & ~x[33] & ~x[34] & ~x[53];
			partial_clause[484] 	= partial_clause_prev[484] & 1'b1;
			partial_clause[485] 	= partial_clause_prev[485] & 1'b1;
			partial_clause[486] 	= partial_clause_prev[486] & ~x[4] & ~x[5] & ~x[17] & ~x[21] & ~x[24] & ~x[26] & ~x[27] & ~x[28] & ~x[39] & ~x[40] & ~x[42] & ~x[51] & ~x[58] & ~x[61];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[34] & ~x[36] & ~x[37] & ~x[55];
			partial_clause[488] 	= partial_clause_prev[488] & ~x[11];
			partial_clause[489] 	= partial_clause_prev[489] & ~x[9] & ~x[13] & ~x[18] & ~x[50] & ~x[51];
			partial_clause[490] 	= partial_clause_prev[490] & 1'b1;
			partial_clause[491] 	= partial_clause_prev[491] & ~x[52];
			partial_clause[492] 	= partial_clause_prev[492] & ~x[3] & ~x[7] & ~x[16] & ~x[34] & ~x[39] & ~x[42] & ~x[44] & ~x[56] & ~x[62];
			partial_clause[493] 	= partial_clause_prev[493] & ~x[51];
			partial_clause[494] 	= partial_clause_prev[494] & ~x[21] & ~x[46] & ~x[51] & ~x[53];
			partial_clause[495] 	= partial_clause_prev[495] & ~x[1] & ~x[2] & ~x[7] & ~x[8] & ~x[62];
			partial_clause[496] 	= partial_clause_prev[496] & 1'b1;
			partial_clause[497] 	= partial_clause_prev[497] & ~x[9];
			partial_clause[498] 	= partial_clause_prev[498] & 1'b1;
			partial_clause[499] 	= partial_clause_prev[499] & ~x[8] & ~x[25] & ~x[59];
		end
	end
endmodule


module HCB_11 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[4] & ~x[6] & ~x[7] & ~x[8] & ~x[10] & ~x[13] & ~x[17] & ~x[19] & ~x[21] & ~x[23] & ~x[29] & ~x[33] & ~x[39] & ~x[43] & ~x[44] & ~x[46] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[59] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[5] & ~x[19] & ~x[34] & ~x[40] & ~x[47];
			partial_clause[2] 	= partial_clause_prev[2] & ~x[45] & ~x[47] & ~x[60];
			partial_clause[3] 	= partial_clause_prev[3] & ~x[33] & ~x[37] & ~x[45] & ~x[46] & ~x[47] & ~x[52] & ~x[53];
			partial_clause[4] 	= partial_clause_prev[4] & ~x[2] & ~x[6] & ~x[11] & ~x[44];
			partial_clause[5] 	= partial_clause_prev[5] & ~x[2] & ~x[4] & ~x[5] & ~x[6] & ~x[9] & ~x[19] & ~x[22] & ~x[32] & ~x[37] & ~x[38] & ~x[50] & ~x[57];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[4] & ~x[8] & ~x[10] & ~x[11] & ~x[12] & ~x[16] & ~x[18] & ~x[32] & ~x[37] & ~x[52] & ~x[56];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[0] & ~x[2] & ~x[5] & ~x[12] & ~x[31] & ~x[44] & ~x[47] & ~x[58] & ~x[62];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[0] & ~x[10] & ~x[11] & ~x[15] & ~x[21] & ~x[23] & ~x[25] & ~x[31] & ~x[33] & ~x[35] & ~x[38] & ~x[44] & ~x[48] & ~x[49] & ~x[54] & ~x[61];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[1] & ~x[2] & ~x[3] & ~x[15] & ~x[21] & ~x[26] & ~x[28] & ~x[31] & ~x[45] & ~x[46] & ~x[51] & ~x[52] & ~x[58] & ~x[60] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[0] & ~x[16] & ~x[23] & ~x[24] & ~x[40] & ~x[44] & ~x[49] & ~x[50] & ~x[55] & ~x[57];
			partial_clause[11] 	= partial_clause_prev[11] & ~x[10] & ~x[11] & ~x[19] & ~x[20] & ~x[26] & ~x[27] & ~x[28] & ~x[38] & ~x[45] & ~x[49] & ~x[50] & ~x[51] & ~x[56] & ~x[57];
			partial_clause[12] 	= partial_clause_prev[12] & ~x[14] & ~x[21] & ~x[41] & ~x[44] & ~x[51] & ~x[53] & ~x[54] & ~x[55] & ~x[58] & ~x[60];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[1] & ~x[7] & ~x[10] & ~x[12] & ~x[14] & ~x[21] & ~x[35] & ~x[39] & ~x[41] & ~x[44] & ~x[50] & ~x[51] & ~x[52] & ~x[54] & ~x[56];
			partial_clause[14] 	= partial_clause_prev[14] & ~x[19];
			partial_clause[15] 	= partial_clause_prev[15] & 1'b1;
			partial_clause[16] 	= partial_clause_prev[16] & ~x[44] & ~x[45] & ~x[55];
			partial_clause[17] 	= partial_clause_prev[17] & ~x[46];
			partial_clause[18] 	= partial_clause_prev[18] & ~x[9] & ~x[46];
			partial_clause[19] 	= partial_clause_prev[19] & ~x[15] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[23] & ~x[25] & ~x[26] & ~x[29] & ~x[38] & ~x[49] & ~x[59];
			partial_clause[20] 	= partial_clause_prev[20] & ~x[0] & ~x[34] & ~x[39];
			partial_clause[21] 	= partial_clause_prev[21] & ~x[29] & ~x[52] & ~x[58] & ~x[63];
			partial_clause[22] 	= partial_clause_prev[22] & ~x[12] & ~x[13] & ~x[23] & ~x[29] & ~x[34] & ~x[41] & ~x[48];
			partial_clause[23] 	= partial_clause_prev[23] & ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[11] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[17] & ~x[18] & ~x[19] & ~x[20] & ~x[22] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & ~x[28] & ~x[31] & ~x[32] & ~x[33] & ~x[34] & ~x[35] & ~x[37] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[45] & ~x[46] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[58] & ~x[59] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[1] & ~x[2] & ~x[3] & ~x[5] & ~x[8] & ~x[12] & ~x[13] & ~x[14] & ~x[15] & ~x[18] & ~x[20] & ~x[21] & ~x[23] & ~x[24] & ~x[25] & ~x[26] & ~x[28] & ~x[30] & ~x[31] & ~x[34] & ~x[36] & ~x[38] & ~x[39] & ~x[45] & ~x[46] & ~x[47] & ~x[49] & ~x[50] & ~x[54] & ~x[59] & ~x[62];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[3] & ~x[4] & ~x[12] & ~x[14] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[27] & ~x[31] & ~x[37] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[46] & ~x[47] & ~x[48] & ~x[51] & ~x[53] & ~x[54] & ~x[55] & ~x[57] & ~x[61];
			partial_clause[26] 	= partial_clause_prev[26] & 1'b1;
			partial_clause[27] 	= partial_clause_prev[27] & ~x[1] & ~x[11] & ~x[14] & ~x[16] & ~x[22] & ~x[28] & ~x[29] & ~x[37] & ~x[44] & ~x[45] & ~x[51];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[1] & ~x[6] & ~x[16] & ~x[23] & ~x[25] & ~x[40];
			partial_clause[29] 	= partial_clause_prev[29] & ~x[24] & ~x[29] & ~x[33] & ~x[35] & ~x[59] & ~x[61] & ~x[62];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[5] & ~x[8] & ~x[21] & ~x[41] & ~x[42] & ~x[52];
			partial_clause[31] 	= partial_clause_prev[31] & ~x[40] & ~x[45] & ~x[47];
			partial_clause[32] 	= partial_clause_prev[32] & ~x[2] & ~x[44];
			partial_clause[33] 	= partial_clause_prev[33] & 1'b1;
			partial_clause[34] 	= partial_clause_prev[34] & ~x[21] & ~x[22] & ~x[28] & ~x[37] & ~x[38] & ~x[40] & ~x[50] & ~x[54] & ~x[56] & ~x[61] & ~x[62];
			partial_clause[35] 	= partial_clause_prev[35] & ~x[3] & ~x[6] & ~x[15] & ~x[18] & ~x[19] & ~x[30] & ~x[38] & ~x[39] & ~x[45] & ~x[48] & ~x[49] & ~x[51] & ~x[58] & ~x[62];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[4] & ~x[7] & ~x[9] & ~x[20] & ~x[28] & ~x[37] & ~x[39] & ~x[42] & ~x[59];
			partial_clause[37] 	= partial_clause_prev[37] & 1'b1;
			partial_clause[38] 	= partial_clause_prev[38] & ~x[10] & ~x[14] & ~x[18] & ~x[19] & ~x[25] & ~x[26] & ~x[40] & ~x[44] & ~x[45] & ~x[48] & ~x[51] & ~x[52] & ~x[56] & ~x[59] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[39] 	= partial_clause_prev[39] & ~x[61];
			partial_clause[40] 	= partial_clause_prev[40] & ~x[14] & ~x[25] & ~x[39] & ~x[42] & ~x[44] & ~x[51] & ~x[54];
			partial_clause[41] 	= partial_clause_prev[41] & 1'b1;
			partial_clause[42] 	= partial_clause_prev[42] & ~x[16] & ~x[37] & ~x[43] & ~x[63];
			partial_clause[43] 	= partial_clause_prev[43] & ~x[41] & ~x[49] & ~x[50] & ~x[51] & ~x[58] & ~x[63];
			partial_clause[44] 	= partial_clause_prev[44] & ~x[55];
			partial_clause[45] 	= partial_clause_prev[45] & ~x[10] & ~x[35] & ~x[46];
			partial_clause[46] 	= partial_clause_prev[46] & ~x[10] & ~x[11] & ~x[15] & ~x[18] & ~x[19] & ~x[27] & ~x[30] & ~x[41] & ~x[44] & ~x[50] & ~x[51] & ~x[52] & ~x[54] & ~x[55] & ~x[63];
			partial_clause[47] 	= partial_clause_prev[47] & ~x[15] & ~x[24] & ~x[26] & ~x[44] & ~x[61];
			partial_clause[48] 	= partial_clause_prev[48] & 1'b1;
			partial_clause[49] 	= partial_clause_prev[49] & ~x[55];
			partial_clause[50] 	= partial_clause_prev[50] & ~x[31];
			partial_clause[51] 	= partial_clause_prev[51] & 1'b1;
			partial_clause[52] 	= partial_clause_prev[52] & 1'b1;
			partial_clause[53] 	= partial_clause_prev[53] & 1'b1;
			partial_clause[54] 	= partial_clause_prev[54] & 1'b1;
			partial_clause[55] 	= partial_clause_prev[55] & 1'b1;
			partial_clause[56] 	= partial_clause_prev[56] & 1'b1;
			partial_clause[57] 	= partial_clause_prev[57] & ~x[9] & ~x[27] & ~x[34] & ~x[36] & ~x[37] & ~x[39] & ~x[40] & ~x[50] & ~x[54] & ~x[55] & ~x[57] & ~x[58];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[12] & ~x[30] & ~x[39] & ~x[42] & ~x[53];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[0] & ~x[1] & ~x[2] & ~x[25] & ~x[27] & ~x[28] & ~x[30] & ~x[34] & ~x[48] & ~x[49] & ~x[54] & ~x[59];
			partial_clause[60] 	= partial_clause_prev[60] & 1'b1;
			partial_clause[61] 	= partial_clause_prev[61] & ~x[10];
			partial_clause[62] 	= partial_clause_prev[62] & ~x[17] & ~x[19] & ~x[54] & ~x[55];
			partial_clause[63] 	= partial_clause_prev[63] & ~x[15] & ~x[36];
			partial_clause[64] 	= partial_clause_prev[64] & ~x[9] & ~x[46];
			partial_clause[65] 	= partial_clause_prev[65] & ~x[5];
			partial_clause[66] 	= partial_clause_prev[66] & 1'b1;
			partial_clause[67] 	= partial_clause_prev[67] & 1'b1;
			partial_clause[68] 	= partial_clause_prev[68] & ~x[27] & ~x[35];
			partial_clause[69] 	= partial_clause_prev[69] & ~x[15] & ~x[17] & ~x[18] & ~x[19] & ~x[31] & ~x[44] & ~x[48] & ~x[56] & ~x[58];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[7] & ~x[10] & ~x[19] & ~x[30] & ~x[32] & ~x[42] & ~x[48] & ~x[57];
			partial_clause[71] 	= partial_clause_prev[71] & ~x[11] & ~x[16] & ~x[61];
			partial_clause[72] 	= partial_clause_prev[72] & ~x[20] & ~x[38];
			partial_clause[73] 	= partial_clause_prev[73] & ~x[50] & ~x[56];
			partial_clause[74] 	= partial_clause_prev[74] & ~x[3] & ~x[7] & ~x[11] & ~x[20] & ~x[29] & ~x[46] & ~x[47] & ~x[51];
			partial_clause[75] 	= partial_clause_prev[75] & ~x[63];
			partial_clause[76] 	= partial_clause_prev[76] & ~x[13] & ~x[18] & ~x[20] & ~x[24] & ~x[38] & ~x[43] & ~x[46] & ~x[58] & ~x[59] & ~x[62];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[2] & ~x[23];
			partial_clause[78] 	= partial_clause_prev[78] & ~x[30] & ~x[36] & ~x[44];
			partial_clause[79] 	= partial_clause_prev[79] & ~x[14] & ~x[22] & ~x[34] & ~x[47] & ~x[53];
			partial_clause[80] 	= partial_clause_prev[80] & 1'b1;
			partial_clause[81] 	= partial_clause_prev[81] & ~x[39];
			partial_clause[82] 	= partial_clause_prev[82] & ~x[6];
			partial_clause[83] 	= partial_clause_prev[83] & 1'b1;
			partial_clause[84] 	= partial_clause_prev[84] & ~x[12] & ~x[53];
			partial_clause[85] 	= partial_clause_prev[85] & ~x[0] & ~x[16] & ~x[21] & ~x[23] & ~x[30] & ~x[35] & ~x[40] & ~x[54];
			partial_clause[86] 	= partial_clause_prev[86] & ~x[1] & ~x[2] & ~x[4] & ~x[13] & ~x[20] & ~x[39] & ~x[40] & ~x[43] & ~x[49] & ~x[51];
			partial_clause[87] 	= partial_clause_prev[87] & ~x[3] & ~x[31] & ~x[58];
			partial_clause[88] 	= partial_clause_prev[88] & ~x[9] & ~x[16] & ~x[27] & ~x[32] & ~x[34] & ~x[40] & ~x[43] & ~x[48] & ~x[53] & ~x[60];
			partial_clause[89] 	= partial_clause_prev[89] & ~x[20] & ~x[51] & ~x[56];
			partial_clause[90] 	= partial_clause_prev[90] & 1'b1;
			partial_clause[91] 	= partial_clause_prev[91] & ~x[13] & ~x[15] & ~x[24] & ~x[51];
			partial_clause[92] 	= partial_clause_prev[92] & ~x[20];
			partial_clause[93] 	= partial_clause_prev[93] & ~x[1] & ~x[8] & ~x[13] & ~x[15] & ~x[21] & ~x[22] & ~x[23] & ~x[25] & ~x[31] & ~x[32] & ~x[33] & ~x[35] & ~x[36] & ~x[40] & ~x[41] & ~x[42] & ~x[44] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[56] & ~x[58] & ~x[59];
			partial_clause[94] 	= partial_clause_prev[94] & 1'b1;
			partial_clause[95] 	= partial_clause_prev[95] & ~x[4] & ~x[7] & ~x[14] & ~x[16] & ~x[28] & ~x[29] & ~x[31] & ~x[32] & ~x[38] & ~x[41] & ~x[42] & ~x[45] & ~x[48] & ~x[54] & ~x[56];
			partial_clause[96] 	= partial_clause_prev[96] & ~x[1];
			partial_clause[97] 	= partial_clause_prev[97] & ~x[15] & ~x[22] & ~x[25] & ~x[30] & ~x[34] & ~x[37] & ~x[39] & ~x[42] & ~x[51] & ~x[55] & ~x[57] & ~x[59] & ~x[60];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[1] & ~x[13] & ~x[14] & ~x[16] & ~x[17] & ~x[18] & ~x[23] & ~x[25] & ~x[27] & ~x[30] & ~x[33] & ~x[35] & ~x[45] & ~x[49] & ~x[50] & ~x[62] & ~x[63];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[1] & ~x[2] & ~x[13] & ~x[16] & ~x[19] & ~x[23] & ~x[25] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & ~x[37] & ~x[38] & ~x[39] & ~x[41] & ~x[46] & ~x[49] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[55] & ~x[56] & ~x[57] & ~x[58] & ~x[61];
			partial_clause[100] 	= partial_clause_prev[100] & ~x[15] & ~x[54] & ~x[55] & ~x[57] & ~x[62];
			partial_clause[101] 	= partial_clause_prev[101] & ~x[54];
			partial_clause[102] 	= partial_clause_prev[102] & ~x[28];
			partial_clause[103] 	= partial_clause_prev[103] & ~x[1] & ~x[13] & ~x[14] & ~x[17] & ~x[20] & ~x[25] & ~x[27] & ~x[30] & ~x[31] & ~x[33] & ~x[37] & ~x[41] & ~x[45] & ~x[46] & ~x[48] & ~x[49] & ~x[54] & ~x[56] & ~x[59] & ~x[62] & ~x[63];
			partial_clause[104] 	= partial_clause_prev[104] & ~x[13] & ~x[17] & ~x[20] & ~x[25] & ~x[27] & ~x[40] & ~x[56] & ~x[59] & ~x[63];
			partial_clause[105] 	= partial_clause_prev[105] & ~x[2] & ~x[4] & ~x[18] & ~x[21] & ~x[28] & ~x[37] & ~x[46] & ~x[47] & ~x[48] & ~x[49] & ~x[62];
			partial_clause[106] 	= partial_clause_prev[106] & ~x[5] & ~x[12] & ~x[26] & ~x[35] & ~x[47] & ~x[53] & ~x[62];
			partial_clause[107] 	= partial_clause_prev[107] & ~x[0] & ~x[13] & ~x[21] & ~x[29] & ~x[34] & ~x[42] & ~x[45] & ~x[48] & ~x[50] & ~x[52] & ~x[54] & ~x[55] & ~x[57];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[1] & ~x[2] & ~x[3] & ~x[7] & ~x[8] & ~x[14] & ~x[15] & ~x[16] & ~x[18] & ~x[22] & ~x[24] & ~x[26] & ~x[27] & ~x[29] & ~x[34] & ~x[37] & ~x[38] & ~x[39] & ~x[41] & ~x[43] & ~x[48] & ~x[49] & ~x[56] & ~x[58] & ~x[63];
			partial_clause[109] 	= partial_clause_prev[109] & 1'b1;
			partial_clause[110] 	= partial_clause_prev[110] & ~x[8] & ~x[37];
			partial_clause[111] 	= partial_clause_prev[111] & 1'b1;
			partial_clause[112] 	= partial_clause_prev[112] & ~x[14] & ~x[25] & ~x[40] & ~x[48] & ~x[51] & ~x[53] & ~x[54];
			partial_clause[113] 	= partial_clause_prev[113] & ~x[6] & ~x[27] & ~x[28] & ~x[36] & ~x[46] & ~x[50] & ~x[58] & ~x[62];
			partial_clause[114] 	= partial_clause_prev[114] & 1'b1;
			partial_clause[115] 	= partial_clause_prev[115] & ~x[21] & ~x[22] & ~x[25] & ~x[26] & ~x[33] & ~x[40] & ~x[45] & ~x[48] & ~x[50] & ~x[55] & ~x[56] & ~x[57];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[14] & ~x[15] & ~x[17] & ~x[26] & ~x[43] & ~x[46] & ~x[47] & ~x[48] & ~x[49] & ~x[53] & ~x[57] & ~x[60];
			partial_clause[117] 	= partial_clause_prev[117] & 1'b1;
			partial_clause[118] 	= partial_clause_prev[118] & ~x[0] & ~x[23] & ~x[43] & ~x[45];
			partial_clause[119] 	= partial_clause_prev[119] & ~x[13] & ~x[15] & ~x[26] & ~x[30] & ~x[36] & ~x[52] & ~x[55] & ~x[62];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[7] & ~x[18] & ~x[20] & ~x[23] & ~x[26] & ~x[29] & ~x[39] & ~x[40] & ~x[45] & ~x[49] & ~x[51] & ~x[52] & ~x[54] & ~x[58] & ~x[59] & ~x[60];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[0] & ~x[8] & ~x[12] & ~x[13] & ~x[14] & ~x[16] & ~x[28] & ~x[31] & ~x[42] & ~x[43] & ~x[52] & ~x[55];
			partial_clause[122] 	= partial_clause_prev[122] & ~x[2] & ~x[18] & ~x[24] & ~x[30] & ~x[38];
			partial_clause[123] 	= partial_clause_prev[123] & ~x[2] & ~x[11] & ~x[13] & ~x[14] & ~x[16] & ~x[17] & ~x[21] & ~x[23] & ~x[24] & ~x[28] & ~x[34] & ~x[43] & ~x[47] & ~x[49] & ~x[51] & ~x[52] & ~x[53] & ~x[57] & ~x[62];
			partial_clause[124] 	= partial_clause_prev[124] & 1'b1;
			partial_clause[125] 	= partial_clause_prev[125] & ~x[0] & ~x[2] & ~x[3] & ~x[8] & ~x[11] & ~x[22] & ~x[26] & ~x[39] & ~x[40];
			partial_clause[126] 	= partial_clause_prev[126] & ~x[10] & ~x[17] & ~x[18] & ~x[25] & ~x[30] & ~x[32] & ~x[35] & ~x[40] & ~x[46] & ~x[48];
			partial_clause[127] 	= partial_clause_prev[127] & ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[6] & ~x[8] & ~x[15] & ~x[16] & ~x[18] & ~x[19] & ~x[21] & ~x[25] & ~x[29] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[42] & ~x[45] & ~x[46] & ~x[48] & ~x[49] & ~x[51] & ~x[61] & ~x[63];
			partial_clause[128] 	= partial_clause_prev[128] & ~x[32];
			partial_clause[129] 	= partial_clause_prev[129] & ~x[7] & ~x[8] & ~x[14] & ~x[15] & ~x[17] & ~x[18] & ~x[22] & ~x[26] & ~x[27] & ~x[29] & ~x[33] & ~x[44] & ~x[45] & ~x[47] & ~x[53] & ~x[57] & ~x[59] & ~x[60];
			partial_clause[130] 	= partial_clause_prev[130] & ~x[2] & ~x[17] & ~x[20] & ~x[26] & ~x[40] & ~x[41] & ~x[45];
			partial_clause[131] 	= partial_clause_prev[131] & 1'b1;
			partial_clause[132] 	= partial_clause_prev[132] & ~x[1] & ~x[8] & ~x[17] & ~x[20] & ~x[21] & ~x[37] & ~x[42] & ~x[46];
			partial_clause[133] 	= partial_clause_prev[133] & ~x[45] & ~x[54];
			partial_clause[134] 	= partial_clause_prev[134] & ~x[14] & ~x[16] & ~x[22] & ~x[23] & ~x[24] & ~x[25] & ~x[28] & ~x[29] & ~x[34] & ~x[35] & ~x[36] & ~x[37] & ~x[38] & ~x[43] & ~x[50] & ~x[54] & ~x[55] & ~x[60] & ~x[63];
			partial_clause[135] 	= partial_clause_prev[135] & ~x[9] & ~x[17] & ~x[23] & ~x[24] & ~x[29] & ~x[62];
			partial_clause[136] 	= partial_clause_prev[136] & ~x[13] & ~x[14] & ~x[15] & ~x[16] & ~x[23] & ~x[32] & ~x[36] & ~x[39] & ~x[52] & ~x[57] & ~x[58];
			partial_clause[137] 	= partial_clause_prev[137] & 1'b1;
			partial_clause[138] 	= partial_clause_prev[138] & 1'b1;
			partial_clause[139] 	= partial_clause_prev[139] & ~x[20] & ~x[23] & ~x[35] & ~x[38] & ~x[39] & ~x[41] & ~x[43] & ~x[45] & ~x[50] & ~x[60] & ~x[63];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[0] & ~x[13] & ~x[16] & ~x[20] & ~x[21] & ~x[23] & ~x[32] & ~x[33] & ~x[34] & ~x[38] & ~x[46] & ~x[52] & ~x[58] & ~x[59] & ~x[61] & ~x[62];
			partial_clause[141] 	= partial_clause_prev[141] & ~x[7] & ~x[10] & ~x[20] & ~x[36] & ~x[38] & ~x[42] & ~x[43] & ~x[47];
			partial_clause[142] 	= partial_clause_prev[142] & ~x[15] & ~x[21] & ~x[22] & ~x[30] & ~x[38] & ~x[39] & ~x[43] & ~x[48] & ~x[54] & ~x[62];
			partial_clause[143] 	= partial_clause_prev[143] & ~x[31] & ~x[41] & ~x[63];
			partial_clause[144] 	= partial_clause_prev[144] & ~x[0] & ~x[23] & ~x[30] & ~x[39] & ~x[40] & ~x[42] & ~x[50] & ~x[53];
			partial_clause[145] 	= partial_clause_prev[145] & ~x[50];
			partial_clause[146] 	= partial_clause_prev[146] & ~x[1] & ~x[7] & ~x[13] & ~x[15] & ~x[17] & ~x[24] & ~x[25] & ~x[28] & ~x[35] & ~x[45] & ~x[58] & ~x[62];
			partial_clause[147] 	= partial_clause_prev[147] & ~x[9] & ~x[21] & ~x[22] & ~x[27] & ~x[36] & ~x[38];
			partial_clause[148] 	= partial_clause_prev[148] & ~x[5] & ~x[19] & ~x[22] & ~x[34] & ~x[36] & ~x[37] & ~x[45] & ~x[47] & ~x[53] & ~x[56] & ~x[61] & ~x[63];
			partial_clause[149] 	= partial_clause_prev[149] & ~x[4] & ~x[7] & ~x[10] & ~x[16] & ~x[20] & ~x[25];
			partial_clause[150] 	= partial_clause_prev[150] & ~x[13] & ~x[17] & ~x[37] & ~x[40] & ~x[44] & ~x[47] & ~x[49] & ~x[50];
			partial_clause[151] 	= partial_clause_prev[151] & 1'b1;
			partial_clause[152] 	= partial_clause_prev[152] & ~x[17] & ~x[21];
			partial_clause[153] 	= partial_clause_prev[153] & ~x[2] & ~x[19] & ~x[35] & ~x[36] & ~x[50] & ~x[55];
			partial_clause[154] 	= partial_clause_prev[154] & ~x[37] & ~x[46] & ~x[62];
			partial_clause[155] 	= partial_clause_prev[155] & 1'b1;
			partial_clause[156] 	= partial_clause_prev[156] & ~x[61];
			partial_clause[157] 	= partial_clause_prev[157] & 1'b1;
			partial_clause[158] 	= partial_clause_prev[158] & ~x[0] & ~x[14] & ~x[16] & ~x[17] & ~x[18] & ~x[22] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & ~x[29] & ~x[41] & ~x[44] & ~x[46] & ~x[47] & ~x[50] & ~x[58];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[0] & ~x[11] & ~x[14] & ~x[15] & ~x[17] & ~x[22] & ~x[24] & ~x[35] & ~x[36] & ~x[37] & ~x[43] & ~x[47] & ~x[53] & ~x[58] & ~x[59] & ~x[60];
			partial_clause[160] 	= partial_clause_prev[160] & ~x[7] & ~x[20] & ~x[46];
			partial_clause[161] 	= partial_clause_prev[161] & ~x[21] & ~x[29] & ~x[30] & ~x[33] & ~x[42] & ~x[59];
			partial_clause[162] 	= partial_clause_prev[162] & ~x[25] & ~x[29] & ~x[35] & ~x[45] & ~x[61];
			partial_clause[163] 	= partial_clause_prev[163] & ~x[3];
			partial_clause[164] 	= partial_clause_prev[164] & ~x[0] & ~x[13] & ~x[28] & ~x[54];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[27] & ~x[41] & ~x[44] & ~x[53];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[4] & ~x[11] & ~x[13] & ~x[16] & ~x[18] & ~x[26] & ~x[27] & ~x[29] & ~x[30] & ~x[32] & ~x[40] & ~x[47] & ~x[52] & ~x[57];
			partial_clause[167] 	= partial_clause_prev[167] & ~x[45] & ~x[56] & ~x[62];
			partial_clause[168] 	= partial_clause_prev[168] & ~x[19] & ~x[25] & ~x[30];
			partial_clause[169] 	= partial_clause_prev[169] & ~x[23];
			partial_clause[170] 	= partial_clause_prev[170] & 1'b1;
			partial_clause[171] 	= partial_clause_prev[171] & ~x[1] & ~x[19] & ~x[22] & ~x[53];
			partial_clause[172] 	= partial_clause_prev[172] & 1'b1;
			partial_clause[173] 	= partial_clause_prev[173] & ~x[16] & ~x[42] & ~x[45] & ~x[52] & ~x[54] & ~x[55] & ~x[58] & ~x[59];
			partial_clause[174] 	= partial_clause_prev[174] & ~x[13] & ~x[16] & ~x[19] & ~x[33] & ~x[48] & ~x[59];
			partial_clause[175] 	= partial_clause_prev[175] & 1'b1;
			partial_clause[176] 	= partial_clause_prev[176] & ~x[32] & ~x[38] & ~x[56];
			partial_clause[177] 	= partial_clause_prev[177] & ~x[14] & ~x[30] & ~x[44] & ~x[55];
			partial_clause[178] 	= partial_clause_prev[178] & ~x[17] & ~x[47] & ~x[57];
			partial_clause[179] 	= partial_clause_prev[179] & 1'b1;
			partial_clause[180] 	= partial_clause_prev[180] & 1'b1;
			partial_clause[181] 	= partial_clause_prev[181] & 1'b1;
			partial_clause[182] 	= partial_clause_prev[182] & 1'b1;
			partial_clause[183] 	= partial_clause_prev[183] & ~x[0] & ~x[2] & ~x[22] & ~x[24] & ~x[28] & ~x[29] & ~x[30] & ~x[45] & ~x[50] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[10] & ~x[18] & ~x[20] & ~x[23] & ~x[25] & ~x[26] & ~x[31] & ~x[34] & ~x[44];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[14] & ~x[18] & ~x[33] & ~x[35] & ~x[40] & ~x[45];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[0] & ~x[5] & ~x[9] & ~x[14] & ~x[20] & ~x[21] & ~x[28] & ~x[31] & ~x[32] & ~x[33] & ~x[35] & ~x[43] & ~x[44] & ~x[45] & ~x[48] & ~x[50] & ~x[61] & ~x[63];
			partial_clause[187] 	= partial_clause_prev[187] & ~x[26] & ~x[55] & ~x[58];
			partial_clause[188] 	= partial_clause_prev[188] & ~x[17] & ~x[55];
			partial_clause[189] 	= partial_clause_prev[189] & 1'b1;
			partial_clause[190] 	= partial_clause_prev[190] & ~x[17] & ~x[23] & ~x[26] & ~x[47];
			partial_clause[191] 	= partial_clause_prev[191] & ~x[11] & ~x[12] & ~x[18] & ~x[19] & ~x[25] & ~x[32] & ~x[42];
			partial_clause[192] 	= partial_clause_prev[192] & ~x[0] & ~x[29] & ~x[30] & ~x[41] & ~x[43];
			partial_clause[193] 	= partial_clause_prev[193] & ~x[3] & ~x[19] & ~x[21] & ~x[24] & ~x[25] & ~x[32];
			partial_clause[194] 	= partial_clause_prev[194] & ~x[5] & ~x[15];
			partial_clause[195] 	= partial_clause_prev[195] & ~x[12] & ~x[19] & ~x[20] & ~x[23] & ~x[26] & ~x[43] & ~x[46] & ~x[47] & ~x[48] & ~x[59] & ~x[61];
			partial_clause[196] 	= partial_clause_prev[196] & ~x[47] & ~x[50] & ~x[59];
			partial_clause[197] 	= partial_clause_prev[197] & ~x[2] & ~x[8] & ~x[9] & ~x[10] & ~x[12] & ~x[13] & ~x[19] & ~x[20] & ~x[24] & ~x[30] & ~x[31] & ~x[33] & ~x[37] & ~x[38] & ~x[39] & ~x[42] & ~x[43] & ~x[45] & ~x[49] & ~x[53] & ~x[63];
			partial_clause[198] 	= partial_clause_prev[198] & 1'b1;
			partial_clause[199] 	= partial_clause_prev[199] & 1'b1;
			partial_clause[200] 	= partial_clause_prev[200] & ~x[38];
			partial_clause[201] 	= partial_clause_prev[201] & ~x[14] & ~x[27] & ~x[28] & ~x[32] & ~x[34] & ~x[39] & ~x[46] & ~x[48] & ~x[53] & ~x[63];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[5] & ~x[7] & ~x[14] & ~x[17] & ~x[20] & ~x[26] & ~x[29] & ~x[30] & ~x[32] & ~x[34] & ~x[35] & ~x[36] & ~x[39] & ~x[41] & ~x[42] & ~x[43] & ~x[54] & ~x[55] & ~x[56] & ~x[58] & ~x[59] & ~x[60] & ~x[63];
			partial_clause[203] 	= partial_clause_prev[203] & ~x[56];
			partial_clause[204] 	= partial_clause_prev[204] & ~x[4] & ~x[5] & ~x[17] & ~x[22] & ~x[30] & ~x[33] & ~x[39] & ~x[42] & ~x[49] & ~x[51] & ~x[62] & ~x[63];
			partial_clause[205] 	= partial_clause_prev[205] & 1'b1;
			partial_clause[206] 	= partial_clause_prev[206] & ~x[14] & ~x[16] & ~x[19] & ~x[28] & ~x[29] & ~x[34] & ~x[35] & ~x[39] & ~x[46] & ~x[51] & ~x[55] & ~x[59];
			partial_clause[207] 	= partial_clause_prev[207] & ~x[1] & ~x[4] & ~x[11] & ~x[36] & ~x[62];
			partial_clause[208] 	= partial_clause_prev[208] & ~x[0] & ~x[26] & ~x[30] & ~x[31] & ~x[32] & ~x[40] & ~x[44];
			partial_clause[209] 	= partial_clause_prev[209] & 1'b1;
			partial_clause[210] 	= partial_clause_prev[210] & ~x[19] & ~x[25] & ~x[31] & ~x[35] & ~x[44] & ~x[49] & ~x[51] & ~x[57];
			partial_clause[211] 	= partial_clause_prev[211] & 1'b1;
			partial_clause[212] 	= partial_clause_prev[212] & ~x[1] & ~x[30] & ~x[34] & ~x[35] & ~x[36] & ~x[41] & ~x[47] & ~x[54] & ~x[61] & ~x[63];
			partial_clause[213] 	= partial_clause_prev[213] & 1'b1;
			partial_clause[214] 	= partial_clause_prev[214] & ~x[8];
			partial_clause[215] 	= partial_clause_prev[215] & ~x[23];
			partial_clause[216] 	= partial_clause_prev[216] & ~x[25] & ~x[36] & ~x[51];
			partial_clause[217] 	= partial_clause_prev[217] & ~x[20] & ~x[26] & ~x[32] & ~x[46] & ~x[49] & ~x[53] & ~x[56] & ~x[63];
			partial_clause[218] 	= partial_clause_prev[218] & ~x[18];
			partial_clause[219] 	= partial_clause_prev[219] & ~x[5];
			partial_clause[220] 	= partial_clause_prev[220] & ~x[17] & ~x[20] & ~x[21] & ~x[24] & ~x[44] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[56] & ~x[60] & ~x[62] & ~x[63];
			partial_clause[221] 	= partial_clause_prev[221] & ~x[30] & ~x[54];
			partial_clause[222] 	= partial_clause_prev[222] & ~x[8];
			partial_clause[223] 	= partial_clause_prev[223] & ~x[13] & ~x[44];
			partial_clause[224] 	= partial_clause_prev[224] & ~x[2] & ~x[4] & ~x[13] & ~x[24] & ~x[28] & ~x[29] & ~x[30] & ~x[33] & ~x[42] & ~x[52] & ~x[58] & ~x[59] & ~x[63];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[1] & ~x[17] & ~x[47] & ~x[49];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[4] & ~x[8] & ~x[20] & ~x[21] & ~x[23] & ~x[25] & ~x[26] & ~x[30] & ~x[37] & ~x[41] & ~x[44] & ~x[46] & ~x[53] & ~x[57] & ~x[59] & ~x[63];
			partial_clause[227] 	= partial_clause_prev[227] & ~x[6] & ~x[9] & ~x[40] & ~x[42] & ~x[55];
			partial_clause[228] 	= partial_clause_prev[228] & ~x[6] & ~x[26] & ~x[49] & ~x[53] & ~x[60];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[2] & ~x[15] & ~x[16] & ~x[18] & ~x[19] & ~x[23] & ~x[24] & ~x[29] & ~x[41] & ~x[46] & ~x[54] & ~x[59] & ~x[60];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[2] & ~x[3] & ~x[15] & ~x[19] & ~x[22] & ~x[23] & ~x[31] & ~x[33] & ~x[34] & ~x[36] & ~x[37] & ~x[42] & ~x[44] & ~x[47] & ~x[52] & ~x[55] & ~x[56] & ~x[59] & ~x[63];
			partial_clause[231] 	= partial_clause_prev[231] & ~x[14] & ~x[18] & ~x[19] & ~x[23] & ~x[33] & ~x[52];
			partial_clause[232] 	= partial_clause_prev[232] & 1'b1;
			partial_clause[233] 	= partial_clause_prev[233] & ~x[4] & ~x[44];
			partial_clause[234] 	= partial_clause_prev[234] & ~x[3] & ~x[8] & ~x[10] & ~x[28];
			partial_clause[235] 	= partial_clause_prev[235] & 1'b1;
			partial_clause[236] 	= partial_clause_prev[236] & 1'b1;
			partial_clause[237] 	= partial_clause_prev[237] & 1'b1;
			partial_clause[238] 	= partial_clause_prev[238] & ~x[22] & ~x[36] & ~x[44];
			partial_clause[239] 	= partial_clause_prev[239] & ~x[1] & ~x[43];
			partial_clause[240] 	= partial_clause_prev[240] & ~x[20] & ~x[21] & ~x[23] & ~x[28] & ~x[44] & ~x[47] & ~x[56] & ~x[59];
			partial_clause[241] 	= partial_clause_prev[241] & 1'b1;
			partial_clause[242] 	= partial_clause_prev[242] & ~x[2] & ~x[5] & ~x[6] & ~x[10] & ~x[15] & ~x[16] & ~x[19] & ~x[30] & ~x[31] & ~x[33] & ~x[40] & ~x[45] & ~x[53];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[2] & ~x[5] & ~x[11] & ~x[12] & ~x[14] & ~x[17] & ~x[19] & ~x[20] & ~x[24] & ~x[25] & ~x[29] & ~x[36] & ~x[41] & ~x[55] & ~x[57] & ~x[59];
			partial_clause[244] 	= partial_clause_prev[244] & ~x[15] & ~x[30];
			partial_clause[245] 	= partial_clause_prev[245] & 1'b1;
			partial_clause[246] 	= partial_clause_prev[246] & ~x[41] & ~x[42] & ~x[45];
			partial_clause[247] 	= partial_clause_prev[247] & ~x[0] & ~x[14] & ~x[15] & ~x[17] & ~x[18] & ~x[20] & ~x[21] & ~x[23] & ~x[29] & ~x[32] & ~x[49] & ~x[50] & ~x[51] & ~x[56] & ~x[58] & ~x[61] & ~x[62];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[1] & ~x[3] & ~x[8] & ~x[9] & ~x[21] & ~x[25] & ~x[26] & ~x[33] & ~x[34] & ~x[36] & ~x[38] & ~x[39] & ~x[46] & ~x[47] & ~x[48] & ~x[50] & ~x[52] & ~x[54];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[11] & ~x[60];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[0] & ~x[14] & ~x[15] & ~x[18] & ~x[20] & ~x[21] & ~x[22] & ~x[24] & ~x[27] & ~x[28] & ~x[30] & ~x[40] & ~x[42] & ~x[44] & ~x[45] & ~x[47] & ~x[48] & ~x[52] & ~x[53] & ~x[54] & ~x[56] & ~x[57] & ~x[58] & ~x[60] & ~x[62];
			partial_clause[251] 	= partial_clause_prev[251] & ~x[18];
			partial_clause[252] 	= partial_clause_prev[252] & ~x[0] & ~x[4] & ~x[6] & ~x[17] & ~x[19] & ~x[25] & ~x[28] & ~x[29] & ~x[31] & ~x[32] & ~x[35] & ~x[38] & ~x[39] & ~x[44] & ~x[48] & ~x[52] & ~x[53] & ~x[55] & ~x[59] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[253] 	= partial_clause_prev[253] & ~x[27] & ~x[61];
			partial_clause[254] 	= partial_clause_prev[254] & ~x[3] & ~x[6] & ~x[17] & ~x[18] & ~x[20] & ~x[29] & ~x[43] & ~x[45] & ~x[49];
			partial_clause[255] 	= partial_clause_prev[255] & ~x[6] & ~x[7] & ~x[11] & ~x[13] & ~x[16] & ~x[22] & ~x[35] & ~x[37] & ~x[44] & ~x[57] & ~x[61];
			partial_clause[256] 	= partial_clause_prev[256] & ~x[43];
			partial_clause[257] 	= partial_clause_prev[257] & ~x[53] & ~x[54] & ~x[55];
			partial_clause[258] 	= partial_clause_prev[258] & ~x[1] & ~x[2] & ~x[18] & ~x[19] & ~x[22] & ~x[25] & ~x[47];
			partial_clause[259] 	= partial_clause_prev[259] & 1'b1;
			partial_clause[260] 	= partial_clause_prev[260] & ~x[1] & ~x[39] & ~x[41] & ~x[58] & ~x[62];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[0] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[15] & ~x[25] & ~x[27] & ~x[29] & ~x[30] & ~x[31];
			partial_clause[262] 	= partial_clause_prev[262] & ~x[18] & ~x[56];
			partial_clause[263] 	= partial_clause_prev[263] & ~x[51] & ~x[59] & ~x[62];
			partial_clause[264] 	= partial_clause_prev[264] & ~x[39];
			partial_clause[265] 	= partial_clause_prev[265] & ~x[27];
			partial_clause[266] 	= partial_clause_prev[266] & ~x[8] & ~x[15] & ~x[23] & ~x[43] & ~x[44] & ~x[50] & ~x[53] & ~x[56];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[1] & ~x[14] & ~x[15] & ~x[19] & ~x[27] & ~x[30] & ~x[36] & ~x[41] & ~x[43] & ~x[44] & ~x[46] & ~x[57];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[1] & ~x[3] & ~x[27] & ~x[28] & ~x[35] & ~x[38] & ~x[39] & ~x[40] & ~x[45] & ~x[47] & ~x[48] & ~x[54] & ~x[55] & ~x[57];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[1] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[10] & ~x[12] & ~x[14] & ~x[16] & ~x[18] & ~x[19] & ~x[20] & ~x[21] & ~x[24] & ~x[33] & ~x[34] & ~x[35] & ~x[37] & ~x[39] & ~x[43] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[52] & ~x[54] & ~x[55] & ~x[57] & ~x[58] & ~x[59] & ~x[60] & ~x[63];
			partial_clause[270] 	= partial_clause_prev[270] & 1'b1;
			partial_clause[271] 	= partial_clause_prev[271] & ~x[3] & ~x[29];
			partial_clause[272] 	= partial_clause_prev[272] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[17] & ~x[26] & ~x[28] & ~x[29] & ~x[33] & ~x[43] & ~x[50] & ~x[51] & ~x[55] & ~x[61] & ~x[63];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[1] & ~x[2] & ~x[5] & ~x[6] & ~x[7] & ~x[11] & ~x[12] & ~x[22] & ~x[24] & ~x[25] & ~x[26] & ~x[27] & ~x[31] & ~x[32] & ~x[33] & ~x[36] & ~x[40] & ~x[43] & ~x[45] & ~x[46] & ~x[47] & ~x[52] & ~x[56] & ~x[57];
			partial_clause[274] 	= partial_clause_prev[274] & ~x[8] & ~x[11] & ~x[22] & ~x[24] & ~x[49] & ~x[55] & ~x[63];
			partial_clause[275] 	= partial_clause_prev[275] & ~x[3] & ~x[4] & ~x[32] & ~x[56] & ~x[57];
			partial_clause[276] 	= partial_clause_prev[276] & ~x[11] & ~x[13] & ~x[33] & ~x[34];
			partial_clause[277] 	= partial_clause_prev[277] & ~x[11] & ~x[22] & ~x[32] & ~x[44];
			partial_clause[278] 	= partial_clause_prev[278] & 1'b1;
			partial_clause[279] 	= partial_clause_prev[279] & ~x[4] & ~x[8] & ~x[17] & ~x[19] & ~x[20] & ~x[21] & ~x[23] & ~x[25] & ~x[32] & ~x[46] & ~x[48] & ~x[49] & ~x[52] & ~x[57] & ~x[62] & ~x[63];
			partial_clause[280] 	= partial_clause_prev[280] & 1'b1;
			partial_clause[281] 	= partial_clause_prev[281] & ~x[0] & ~x[4] & ~x[5] & ~x[16] & ~x[17] & ~x[18] & ~x[23] & ~x[31] & ~x[43] & ~x[46] & ~x[54];
			partial_clause[282] 	= partial_clause_prev[282] & ~x[0] & ~x[2] & ~x[4] & ~x[16] & ~x[57];
			partial_clause[283] 	= partial_clause_prev[283] & ~x[15] & ~x[59];
			partial_clause[284] 	= partial_clause_prev[284] & ~x[43];
			partial_clause[285] 	= partial_clause_prev[285] & 1'b1;
			partial_clause[286] 	= partial_clause_prev[286] & ~x[54];
			partial_clause[287] 	= partial_clause_prev[287] & ~x[1] & ~x[2] & ~x[14] & ~x[16] & ~x[19] & ~x[23] & ~x[26] & ~x[28] & ~x[34] & ~x[35] & ~x[40] & ~x[45] & ~x[50] & ~x[52] & ~x[60] & ~x[61];
			partial_clause[288] 	= partial_clause_prev[288] & ~x[19] & ~x[53];
			partial_clause[289] 	= partial_clause_prev[289] & ~x[3] & ~x[43] & ~x[44] & ~x[45] & ~x[56];
			partial_clause[290] 	= partial_clause_prev[290] & ~x[31] & ~x[36] & ~x[37] & ~x[59];
			partial_clause[291] 	= partial_clause_prev[291] & ~x[9] & ~x[53];
			partial_clause[292] 	= partial_clause_prev[292] & ~x[26] & ~x[48] & ~x[53];
			partial_clause[293] 	= partial_clause_prev[293] & ~x[19] & ~x[24] & ~x[39] & ~x[52] & ~x[53] & ~x[59];
			partial_clause[294] 	= partial_clause_prev[294] & ~x[57];
			partial_clause[295] 	= partial_clause_prev[295] & ~x[8] & ~x[10] & ~x[29] & ~x[32] & ~x[45];
			partial_clause[296] 	= partial_clause_prev[296] & ~x[51];
			partial_clause[297] 	= partial_clause_prev[297] & ~x[21] & ~x[25] & ~x[40];
			partial_clause[298] 	= partial_clause_prev[298] & 1'b1;
			partial_clause[299] 	= partial_clause_prev[299] & ~x[1] & ~x[22] & ~x[29] & ~x[33] & ~x[51] & ~x[59];
			partial_clause[300] 	= partial_clause_prev[300] & ~x[0] & ~x[1] & ~x[4] & ~x[5] & ~x[12] & ~x[13] & ~x[25] & ~x[41] & ~x[59];
			partial_clause[301] 	= partial_clause_prev[301] & ~x[27] & ~x[43] & ~x[48] & ~x[54] & ~x[57];
			partial_clause[302] 	= partial_clause_prev[302] & ~x[18] & ~x[36] & ~x[40] & ~x[54] & ~x[62];
			partial_clause[303] 	= partial_clause_prev[303] & ~x[2] & ~x[50];
			partial_clause[304] 	= partial_clause_prev[304] & ~x[1] & ~x[7] & ~x[9] & ~x[32] & ~x[55] & ~x[57] & ~x[63];
			partial_clause[305] 	= partial_clause_prev[305] & ~x[8] & ~x[17] & ~x[21] & ~x[31];
			partial_clause[306] 	= partial_clause_prev[306] & ~x[2] & ~x[14] & ~x[23] & ~x[48] & ~x[49] & ~x[50] & ~x[52];
			partial_clause[307] 	= partial_clause_prev[307] & ~x[4] & ~x[11] & ~x[26] & ~x[27] & ~x[29] & ~x[38] & ~x[46] & ~x[49] & ~x[50] & ~x[63];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[5] & ~x[6] & ~x[19] & ~x[25] & ~x[26] & ~x[28] & ~x[29] & ~x[42] & ~x[43] & ~x[47] & ~x[55];
			partial_clause[309] 	= partial_clause_prev[309] & ~x[2] & ~x[6] & ~x[9] & ~x[11] & ~x[13] & ~x[27] & ~x[31] & ~x[35] & ~x[43] & ~x[57] & ~x[59];
			partial_clause[310] 	= partial_clause_prev[310] & 1'b1;
			partial_clause[311] 	= partial_clause_prev[311] & ~x[11] & ~x[24] & ~x[40] & ~x[43] & ~x[52] & ~x[54];
			partial_clause[312] 	= partial_clause_prev[312] & 1'b1;
			partial_clause[313] 	= partial_clause_prev[313] & ~x[22] & ~x[23] & ~x[28] & ~x[37];
			partial_clause[314] 	= partial_clause_prev[314] & ~x[16] & ~x[28] & ~x[33] & ~x[60];
			partial_clause[315] 	= partial_clause_prev[315] & ~x[24] & ~x[55];
			partial_clause[316] 	= partial_clause_prev[316] & ~x[2] & ~x[5] & ~x[6] & ~x[27] & ~x[30] & ~x[31] & ~x[34] & ~x[35] & ~x[37] & ~x[47] & ~x[56] & ~x[59] & ~x[60];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[1] & ~x[4] & ~x[10] & ~x[11] & ~x[26] & ~x[51] & ~x[53] & ~x[55];
			partial_clause[318] 	= partial_clause_prev[318] & ~x[22];
			partial_clause[319] 	= partial_clause_prev[319] & ~x[31] & ~x[41];
			partial_clause[320] 	= partial_clause_prev[320] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[15] & ~x[17] & ~x[22] & ~x[27] & ~x[31] & ~x[34] & ~x[35] & ~x[45] & ~x[46] & ~x[49] & ~x[50];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[1] & ~x[28] & ~x[37] & ~x[47] & ~x[60] & ~x[61];
			partial_clause[322] 	= partial_clause_prev[322] & ~x[10] & ~x[14] & ~x[16] & ~x[20] & ~x[27] & ~x[29] & ~x[30] & ~x[31] & ~x[44] & ~x[47] & ~x[59];
			partial_clause[323] 	= partial_clause_prev[323] & ~x[20] & ~x[31] & ~x[57];
			partial_clause[324] 	= partial_clause_prev[324] & ~x[11] & ~x[13];
			partial_clause[325] 	= partial_clause_prev[325] & ~x[0] & ~x[4] & ~x[5] & ~x[6] & ~x[9] & ~x[10] & ~x[12] & ~x[15] & ~x[19] & ~x[20] & ~x[28] & ~x[29] & ~x[31] & ~x[32] & ~x[35] & ~x[37] & ~x[39] & ~x[40] & ~x[43] & ~x[48] & ~x[51] & ~x[53] & ~x[54] & ~x[55] & ~x[57] & ~x[58] & ~x[59] & ~x[61] & ~x[62];
			partial_clause[326] 	= partial_clause_prev[326] & ~x[3] & ~x[29] & ~x[31] & ~x[33] & ~x[35] & ~x[47] & ~x[52] & ~x[62];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[6] & ~x[22] & ~x[40] & ~x[45];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[9] & ~x[44] & ~x[62];
			partial_clause[329] 	= partial_clause_prev[329] & 1'b1;
			partial_clause[330] 	= partial_clause_prev[330] & ~x[14] & ~x[36] & ~x[47] & ~x[60] & ~x[61];
			partial_clause[331] 	= partial_clause_prev[331] & ~x[2] & ~x[18] & ~x[21] & ~x[50] & ~x[58];
			partial_clause[332] 	= partial_clause_prev[332] & ~x[4] & ~x[6] & ~x[26] & ~x[30] & ~x[32] & ~x[37] & ~x[49] & ~x[56] & ~x[62] & ~x[63];
			partial_clause[333] 	= partial_clause_prev[333] & ~x[29] & ~x[43] & ~x[63];
			partial_clause[334] 	= partial_clause_prev[334] & ~x[20] & ~x[27] & ~x[34] & ~x[48] & ~x[62];
			partial_clause[335] 	= partial_clause_prev[335] & ~x[30] & ~x[49];
			partial_clause[336] 	= partial_clause_prev[336] & 1'b1;
			partial_clause[337] 	= partial_clause_prev[337] & ~x[3] & ~x[5] & ~x[13] & ~x[14] & ~x[18] & ~x[22] & ~x[25] & ~x[26] & ~x[29] & ~x[37] & ~x[41] & ~x[49] & ~x[55];
			partial_clause[338] 	= partial_clause_prev[338] & 1'b1;
			partial_clause[339] 	= partial_clause_prev[339] & ~x[0] & ~x[4] & ~x[16] & ~x[23] & ~x[26] & ~x[27] & ~x[28] & ~x[31] & ~x[32] & ~x[41] & ~x[45] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[59] & ~x[62];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[18] & ~x[23] & ~x[27] & ~x[47] & ~x[48] & ~x[52] & ~x[56];
			partial_clause[341] 	= partial_clause_prev[341] & 1'b1;
			partial_clause[342] 	= partial_clause_prev[342] & ~x[11] & ~x[12] & ~x[16] & ~x[19] & ~x[23] & ~x[30] & ~x[32] & ~x[34] & ~x[50];
			partial_clause[343] 	= partial_clause_prev[343] & ~x[1] & ~x[25] & ~x[26] & ~x[52] & ~x[58] & ~x[62];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[7] & ~x[9] & ~x[19] & ~x[30] & ~x[35] & ~x[49] & ~x[61];
			partial_clause[345] 	= partial_clause_prev[345] & ~x[9] & ~x[10] & ~x[11] & ~x[22] & ~x[54];
			partial_clause[346] 	= partial_clause_prev[346] & ~x[27] & ~x[50] & ~x[51];
			partial_clause[347] 	= partial_clause_prev[347] & ~x[24] & ~x[31] & ~x[37] & ~x[45] & ~x[48] & ~x[52] & ~x[57] & ~x[60];
			partial_clause[348] 	= partial_clause_prev[348] & ~x[44] & ~x[47] & ~x[55];
			partial_clause[349] 	= partial_clause_prev[349] & ~x[21] & ~x[28] & ~x[29] & ~x[41] & ~x[59];
			partial_clause[350] 	= partial_clause_prev[350] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[20] & ~x[21] & ~x[25] & ~x[27] & ~x[29] & ~x[31] & ~x[32] & ~x[36] & ~x[37] & ~x[40] & ~x[41] & ~x[43] & ~x[44] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[54] & ~x[55] & ~x[56] & ~x[59] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[351] 	= partial_clause_prev[351] & 1'b1;
			partial_clause[352] 	= partial_clause_prev[352] & 1'b1;
			partial_clause[353] 	= partial_clause_prev[353] & ~x[22];
			partial_clause[354] 	= partial_clause_prev[354] & ~x[0] & ~x[1] & ~x[4] & ~x[7] & ~x[10] & ~x[14] & ~x[30] & ~x[34] & ~x[39] & ~x[41] & ~x[46] & ~x[47] & ~x[54];
			partial_clause[355] 	= partial_clause_prev[355] & ~x[6] & ~x[21] & ~x[26] & ~x[27] & ~x[33];
			partial_clause[356] 	= partial_clause_prev[356] & ~x[6] & ~x[11] & ~x[28] & ~x[30] & ~x[34] & ~x[35];
			partial_clause[357] 	= partial_clause_prev[357] & ~x[24];
			partial_clause[358] 	= partial_clause_prev[358] & ~x[7] & ~x[18] & ~x[27] & ~x[39] & ~x[45] & ~x[46] & ~x[57];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[2] & ~x[9] & ~x[17] & ~x[18] & ~x[34] & ~x[36] & ~x[56] & ~x[63];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[2] & ~x[23] & ~x[28] & ~x[48] & ~x[49] & ~x[53] & ~x[54] & ~x[56] & ~x[58] & ~x[61] & ~x[62];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[23] & ~x[24] & ~x[32] & ~x[49] & ~x[59];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[34] & ~x[54] & ~x[57];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[1] & ~x[3] & ~x[7] & ~x[19] & ~x[20] & ~x[22] & ~x[31] & ~x[38] & ~x[41] & ~x[44] & ~x[48] & ~x[52] & ~x[54] & ~x[63];
			partial_clause[364] 	= partial_clause_prev[364] & ~x[11] & ~x[12] & ~x[24] & ~x[26] & ~x[35] & ~x[44] & ~x[48] & ~x[54] & ~x[61];
			partial_clause[365] 	= partial_clause_prev[365] & 1'b1;
			partial_clause[366] 	= partial_clause_prev[366] & ~x[8] & ~x[30] & ~x[40] & ~x[46] & ~x[47] & ~x[52] & ~x[53] & ~x[54] & ~x[58];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[20] & ~x[21] & ~x[25] & ~x[26] & ~x[28] & ~x[44];
			partial_clause[368] 	= partial_clause_prev[368] & 1'b1;
			partial_clause[369] 	= partial_clause_prev[369] & ~x[22] & ~x[24] & ~x[29] & ~x[53];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[3] & ~x[46] & ~x[55] & ~x[62];
			partial_clause[371] 	= partial_clause_prev[371] & ~x[16];
			partial_clause[372] 	= partial_clause_prev[372] & ~x[17] & ~x[30] & ~x[32] & ~x[45] & ~x[57] & ~x[59];
			partial_clause[373] 	= partial_clause_prev[373] & ~x[38];
			partial_clause[374] 	= partial_clause_prev[374] & ~x[49];
			partial_clause[375] 	= partial_clause_prev[375] & 1'b1;
			partial_clause[376] 	= partial_clause_prev[376] & ~x[44] & ~x[51] & ~x[62] & ~x[63];
			partial_clause[377] 	= partial_clause_prev[377] & ~x[1] & ~x[5] & ~x[32];
			partial_clause[378] 	= partial_clause_prev[378] & ~x[1] & ~x[34];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[37] & ~x[46] & ~x[56] & ~x[62];
			partial_clause[380] 	= partial_clause_prev[380] & 1'b1;
			partial_clause[381] 	= partial_clause_prev[381] & ~x[1] & ~x[2] & ~x[6] & ~x[10] & ~x[11] & ~x[13] & ~x[15] & ~x[17] & ~x[20] & ~x[23] & ~x[49] & ~x[54] & ~x[55] & ~x[61] & ~x[62] & ~x[63];
			partial_clause[382] 	= partial_clause_prev[382] & 1'b1;
			partial_clause[383] 	= partial_clause_prev[383] & ~x[62];
			partial_clause[384] 	= partial_clause_prev[384] & 1'b1;
			partial_clause[385] 	= partial_clause_prev[385] & 1'b1;
			partial_clause[386] 	= partial_clause_prev[386] & 1'b1;
			partial_clause[387] 	= partial_clause_prev[387] & ~x[3] & ~x[4] & ~x[6] & ~x[11] & ~x[12] & ~x[14] & ~x[20] & ~x[23] & ~x[24] & ~x[26] & ~x[33] & ~x[36] & ~x[38] & ~x[41] & ~x[42] & ~x[46] & ~x[50] & ~x[53] & ~x[55] & ~x[59];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[0] & ~x[1] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[18] & ~x[19] & ~x[23] & ~x[24] & ~x[29] & ~x[31] & ~x[32] & ~x[34] & ~x[39] & ~x[41] & ~x[43] & ~x[45] & ~x[51] & ~x[54] & ~x[55] & ~x[56] & ~x[60];
			partial_clause[389] 	= partial_clause_prev[389] & 1'b1;
			partial_clause[390] 	= partial_clause_prev[390] & ~x[3] & ~x[6] & ~x[8] & ~x[20] & ~x[24] & ~x[29] & ~x[42] & ~x[50] & ~x[52] & ~x[56] & ~x[63];
			partial_clause[391] 	= partial_clause_prev[391] & 1'b1;
			partial_clause[392] 	= partial_clause_prev[392] & 1'b1;
			partial_clause[393] 	= partial_clause_prev[393] & 1'b1;
			partial_clause[394] 	= partial_clause_prev[394] & ~x[2] & ~x[28] & ~x[45] & ~x[48];
			partial_clause[395] 	= partial_clause_prev[395] & ~x[5] & ~x[8];
			partial_clause[396] 	= partial_clause_prev[396] & ~x[30];
			partial_clause[397] 	= partial_clause_prev[397] & ~x[25];
			partial_clause[398] 	= partial_clause_prev[398] & 1'b1;
			partial_clause[399] 	= partial_clause_prev[399] & 1'b1;
			partial_clause[400] 	= partial_clause_prev[400] & ~x[17] & ~x[26] & ~x[28] & ~x[33] & ~x[38] & ~x[41] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[62];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[13] & ~x[17] & ~x[22] & ~x[29] & ~x[31] & ~x[45] & ~x[48] & ~x[55] & ~x[62];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[5] & ~x[13] & ~x[14] & ~x[17] & ~x[20] & ~x[22] & ~x[23] & ~x[29] & ~x[34] & ~x[40] & ~x[43] & ~x[49] & ~x[58] & ~x[63];
			partial_clause[403] 	= partial_clause_prev[403] & ~x[31] & ~x[57];
			partial_clause[404] 	= partial_clause_prev[404] & 1'b1;
			partial_clause[405] 	= partial_clause_prev[405] & ~x[16] & ~x[21] & ~x[25] & ~x[29] & ~x[54];
			partial_clause[406] 	= partial_clause_prev[406] & ~x[34] & ~x[35] & ~x[37] & ~x[51];
			partial_clause[407] 	= partial_clause_prev[407] & ~x[18] & ~x[25];
			partial_clause[408] 	= partial_clause_prev[408] & ~x[20] & ~x[27] & ~x[40];
			partial_clause[409] 	= partial_clause_prev[409] & ~x[0] & ~x[1] & ~x[4] & ~x[6] & ~x[14] & ~x[15] & ~x[18] & ~x[20] & ~x[23] & ~x[26] & ~x[31] & ~x[33] & ~x[36] & ~x[37] & ~x[38] & ~x[40] & ~x[43] & ~x[52] & ~x[54] & ~x[57] & ~x[59] & ~x[63];
			partial_clause[410] 	= partial_clause_prev[410] & ~x[4] & ~x[6] & ~x[7] & ~x[13] & ~x[14] & ~x[16] & ~x[31] & ~x[37] & ~x[38] & ~x[44];
			partial_clause[411] 	= partial_clause_prev[411] & ~x[2] & ~x[6] & ~x[42] & ~x[43] & ~x[54] & ~x[56] & ~x[57] & ~x[61];
			partial_clause[412] 	= partial_clause_prev[412] & ~x[3] & ~x[9] & ~x[17] & ~x[19] & ~x[21] & ~x[28] & ~x[30] & ~x[34] & ~x[42] & ~x[45] & ~x[46] & ~x[47] & ~x[48] & ~x[49] & ~x[51] & ~x[53] & ~x[55] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[413] 	= partial_clause_prev[413] & 1'b1;
			partial_clause[414] 	= partial_clause_prev[414] & ~x[0] & ~x[1] & ~x[3] & ~x[7] & ~x[8] & ~x[9] & ~x[11] & ~x[13] & ~x[22] & ~x[24] & ~x[27] & ~x[28] & ~x[33] & ~x[35] & ~x[39] & ~x[42] & ~x[43] & ~x[45] & ~x[61] & ~x[62];
			partial_clause[415] 	= partial_clause_prev[415] & ~x[53] & ~x[62];
			partial_clause[416] 	= partial_clause_prev[416] & ~x[8] & ~x[9] & ~x[10] & ~x[19] & ~x[20] & ~x[25] & ~x[26] & ~x[29] & ~x[30] & ~x[36] & ~x[39] & ~x[46] & ~x[51] & ~x[53] & ~x[54] & ~x[55] & ~x[56] & ~x[57] & ~x[61];
			partial_clause[417] 	= partial_clause_prev[417] & ~x[9] & ~x[12] & ~x[32] & ~x[45] & ~x[47] & ~x[48] & ~x[57] & ~x[60];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[5] & ~x[20] & ~x[23] & ~x[25] & ~x[27] & ~x[29] & ~x[34] & ~x[53] & ~x[56] & ~x[58] & ~x[59] & ~x[60] & ~x[61];
			partial_clause[419] 	= partial_clause_prev[419] & 1'b1;
			partial_clause[420] 	= partial_clause_prev[420] & ~x[39];
			partial_clause[421] 	= partial_clause_prev[421] & ~x[1] & ~x[16] & ~x[24] & ~x[32] & ~x[34] & ~x[47] & ~x[53] & ~x[54] & ~x[55];
			partial_clause[422] 	= partial_clause_prev[422] & ~x[2] & ~x[22] & ~x[43] & ~x[50];
			partial_clause[423] 	= partial_clause_prev[423] & ~x[50] & ~x[51] & ~x[58];
			partial_clause[424] 	= partial_clause_prev[424] & ~x[59];
			partial_clause[425] 	= partial_clause_prev[425] & ~x[9] & ~x[11] & ~x[23] & ~x[45];
			partial_clause[426] 	= partial_clause_prev[426] & ~x[0] & ~x[14] & ~x[18] & ~x[20] & ~x[22] & ~x[23] & ~x[26] & ~x[31] & ~x[46] & ~x[55] & ~x[56] & ~x[60] & ~x[61] & ~x[63];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[20] & ~x[21] & ~x[24] & ~x[26] & ~x[27] & ~x[52] & ~x[53] & ~x[55] & ~x[56] & ~x[57] & ~x[59];
			partial_clause[428] 	= partial_clause_prev[428] & ~x[9] & ~x[45];
			partial_clause[429] 	= partial_clause_prev[429] & 1'b1;
			partial_clause[430] 	= partial_clause_prev[430] & ~x[0] & ~x[4] & ~x[8] & ~x[13] & ~x[17] & ~x[18] & ~x[26] & ~x[27] & ~x[32] & ~x[51] & ~x[56] & ~x[58] & ~x[59] & ~x[60];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[19] & ~x[56] & ~x[58];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[19] & ~x[31] & ~x[32] & ~x[37] & ~x[38] & ~x[52] & ~x[56] & ~x[59];
			partial_clause[433] 	= partial_clause_prev[433] & ~x[20] & ~x[56];
			partial_clause[434] 	= partial_clause_prev[434] & ~x[1] & ~x[55];
			partial_clause[435] 	= partial_clause_prev[435] & ~x[0] & ~x[14] & ~x[15] & ~x[16] & ~x[18] & ~x[19] & ~x[23] & ~x[28] & ~x[31] & ~x[32] & ~x[39] & ~x[43] & ~x[48] & ~x[49] & ~x[50] & ~x[56] & ~x[59] & ~x[61] & ~x[62];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[11] & ~x[12] & ~x[13] & ~x[18] & ~x[19] & ~x[25] & ~x[26] & ~x[44] & ~x[45] & ~x[51];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[1] & ~x[2] & ~x[10] & ~x[14] & ~x[21] & ~x[23] & ~x[25] & ~x[34] & ~x[40] & ~x[41] & ~x[42] & ~x[45] & ~x[48] & ~x[52] & ~x[60] & ~x[62];
			partial_clause[438] 	= partial_clause_prev[438] & 1'b1;
			partial_clause[439] 	= partial_clause_prev[439] & ~x[1] & ~x[4] & ~x[42] & ~x[45];
			partial_clause[440] 	= partial_clause_prev[440] & 1'b1;
			partial_clause[441] 	= partial_clause_prev[441] & ~x[5] & ~x[54] & ~x[63];
			partial_clause[442] 	= partial_clause_prev[442] & 1'b1;
			partial_clause[443] 	= partial_clause_prev[443] & ~x[19] & ~x[21] & ~x[22] & ~x[25] & ~x[46] & ~x[47] & ~x[52];
			partial_clause[444] 	= partial_clause_prev[444] & 1'b1;
			partial_clause[445] 	= partial_clause_prev[445] & ~x[18];
			partial_clause[446] 	= partial_clause_prev[446] & ~x[2] & ~x[26] & ~x[36] & ~x[44] & ~x[45];
			partial_clause[447] 	= partial_clause_prev[447] & ~x[0] & ~x[15] & ~x[19] & ~x[27] & ~x[35] & ~x[42] & ~x[54] & ~x[62];
			partial_clause[448] 	= partial_clause_prev[448] & 1'b1;
			partial_clause[449] 	= partial_clause_prev[449] & ~x[6] & ~x[26] & ~x[39] & ~x[41] & ~x[51];
			partial_clause[450] 	= partial_clause_prev[450] & ~x[10] & ~x[32] & ~x[51] & ~x[62];
			partial_clause[451] 	= partial_clause_prev[451] & 1'b1;
			partial_clause[452] 	= partial_clause_prev[452] & 1'b1;
			partial_clause[453] 	= partial_clause_prev[453] & ~x[33] & ~x[35];
			partial_clause[454] 	= partial_clause_prev[454] & ~x[13] & ~x[14] & ~x[21] & ~x[23] & ~x[56];
			partial_clause[455] 	= partial_clause_prev[455] & ~x[15] & ~x[23] & ~x[40] & ~x[42] & ~x[48] & ~x[57];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[2] & ~x[11] & ~x[18] & ~x[22] & ~x[38] & ~x[39] & ~x[43] & ~x[45] & ~x[46] & ~x[54];
			partial_clause[457] 	= partial_clause_prev[457] & ~x[42];
			partial_clause[458] 	= partial_clause_prev[458] & ~x[15] & ~x[22] & ~x[27] & ~x[37] & ~x[41] & ~x[46] & ~x[47] & ~x[51] & ~x[52] & ~x[62] & ~x[63];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[14] & ~x[16] & ~x[34] & ~x[36] & ~x[41] & ~x[45] & ~x[48] & ~x[51] & ~x[59];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[2] & ~x[5] & ~x[7] & ~x[8] & ~x[18] & ~x[24] & ~x[25] & ~x[29] & ~x[30] & ~x[37] & ~x[38] & ~x[43] & ~x[53] & ~x[55] & ~x[59];
			partial_clause[461] 	= partial_clause_prev[461] & ~x[58] & ~x[59] & ~x[62];
			partial_clause[462] 	= partial_clause_prev[462] & ~x[39] & ~x[62];
			partial_clause[463] 	= partial_clause_prev[463] & 1'b1;
			partial_clause[464] 	= partial_clause_prev[464] & ~x[3] & ~x[4] & ~x[16] & ~x[20] & ~x[22] & ~x[44] & ~x[51] & ~x[52] & ~x[54];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[3] & ~x[6] & ~x[31] & ~x[34] & ~x[35] & ~x[40] & ~x[41] & ~x[48] & ~x[50] & ~x[52] & ~x[56] & ~x[57] & ~x[60] & ~x[63];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[1] & ~x[2] & ~x[4] & ~x[9] & ~x[23] & ~x[25] & ~x[27] & ~x[29] & ~x[34] & ~x[35] & ~x[37] & ~x[40] & ~x[42] & ~x[45] & ~x[55] & ~x[59] & ~x[60];
			partial_clause[467] 	= partial_clause_prev[467] & ~x[7] & ~x[50] & ~x[58];
			partial_clause[468] 	= partial_clause_prev[468] & ~x[15] & ~x[28] & ~x[39] & ~x[50];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[2] & ~x[24] & ~x[44] & ~x[52];
			partial_clause[470] 	= partial_clause_prev[470] & ~x[49];
			partial_clause[471] 	= partial_clause_prev[471] & ~x[4] & ~x[7] & ~x[10] & ~x[13] & ~x[17] & ~x[18] & ~x[20] & ~x[22] & ~x[23] & ~x[26] & ~x[41] & ~x[47] & ~x[48] & ~x[49] & ~x[60] & ~x[62];
			partial_clause[472] 	= partial_clause_prev[472] & ~x[55];
			partial_clause[473] 	= partial_clause_prev[473] & ~x[4] & ~x[14] & ~x[15] & ~x[17] & ~x[22] & ~x[26] & ~x[32] & ~x[41] & ~x[42] & ~x[46] & ~x[50] & ~x[51] & ~x[56];
			partial_clause[474] 	= partial_clause_prev[474] & ~x[19] & ~x[31];
			partial_clause[475] 	= partial_clause_prev[475] & ~x[18] & ~x[59];
			partial_clause[476] 	= partial_clause_prev[476] & 1'b1;
			partial_clause[477] 	= partial_clause_prev[477] & ~x[3] & ~x[20] & ~x[31] & ~x[41] & ~x[51] & ~x[52] & ~x[55] & ~x[63];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[4] & ~x[13] & ~x[14] & ~x[23] & ~x[25] & ~x[27] & ~x[29] & ~x[33] & ~x[35] & ~x[38] & ~x[43] & ~x[51] & ~x[52] & ~x[54] & ~x[56] & ~x[61];
			partial_clause[479] 	= partial_clause_prev[479] & ~x[49];
			partial_clause[480] 	= partial_clause_prev[480] & ~x[0] & ~x[1] & ~x[3] & ~x[4] & ~x[14] & ~x[15] & ~x[17] & ~x[19] & ~x[20] & ~x[21] & ~x[22] & ~x[23] & ~x[25] & ~x[26] & ~x[27] & ~x[28] & ~x[29] & ~x[30] & ~x[31] & ~x[32] & ~x[33] & ~x[35] & ~x[37] & ~x[38] & ~x[39] & ~x[40] & ~x[41] & ~x[42] & ~x[43] & ~x[44] & ~x[45] & ~x[46] & ~x[47] & ~x[48] & ~x[49] & ~x[50] & ~x[51] & ~x[52] & ~x[53] & ~x[54] & ~x[57] & ~x[58] & ~x[59] & ~x[60] & ~x[61] & ~x[62];
			partial_clause[481] 	= partial_clause_prev[481] & ~x[3] & ~x[20] & ~x[37] & ~x[40];
			partial_clause[482] 	= partial_clause_prev[482] & ~x[2] & ~x[4] & ~x[44] & ~x[49];
			partial_clause[483] 	= partial_clause_prev[483] & ~x[33] & ~x[35] & ~x[36] & ~x[58];
			partial_clause[484] 	= partial_clause_prev[484] & ~x[2] & ~x[7] & ~x[19] & ~x[30] & ~x[37] & ~x[63];
			partial_clause[485] 	= partial_clause_prev[485] & ~x[63];
			partial_clause[486] 	= partial_clause_prev[486] & ~x[0] & ~x[1] & ~x[2] & ~x[9] & ~x[11] & ~x[14] & ~x[15] & ~x[21] & ~x[25] & ~x[31] & ~x[32] & ~x[34] & ~x[42] & ~x[58] & ~x[62];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[11] & ~x[16] & ~x[24] & ~x[28] & ~x[32] & ~x[40] & ~x[56];
			partial_clause[488] 	= partial_clause_prev[488] & ~x[5];
			partial_clause[489] 	= partial_clause_prev[489] & ~x[10];
			partial_clause[490] 	= partial_clause_prev[490] & 1'b1;
			partial_clause[491] 	= partial_clause_prev[491] & ~x[0] & ~x[46];
			partial_clause[492] 	= partial_clause_prev[492] & ~x[9] & ~x[13] & ~x[25] & ~x[27] & ~x[28] & ~x[46] & ~x[61];
			partial_clause[493] 	= partial_clause_prev[493] & ~x[57] & ~x[63];
			partial_clause[494] 	= partial_clause_prev[494] & ~x[18];
			partial_clause[495] 	= partial_clause_prev[495] & ~x[29] & ~x[30] & ~x[32] & ~x[37] & ~x[47] & ~x[48] & ~x[63];
			partial_clause[496] 	= partial_clause_prev[496] & 1'b1;
			partial_clause[497] 	= partial_clause_prev[497] & 1'b1;
			partial_clause[498] 	= partial_clause_prev[498] & 1'b1;
			partial_clause[499] 	= partial_clause_prev[499] & ~x[13] & ~x[15] & ~x[27] & ~x[43] & ~x[48] & ~x[51];
		end
	end
endmodule


module HCB_12 (x, partial_clause, partial_clause_prev, clk, valid);
	input	logic [499:0] partial_clause_prev;
	output	logic[499:0] partial_clause;
	input	logic clk;
	input	logic [63:0] x;
	input	logic valid;
	always @(posedge clk) begin
		if(valid) begin
			partial_clause[0] 	= partial_clause_prev[0] & ~x[0] & ~x[7] & ~x[15];
			partial_clause[1] 	= partial_clause_prev[1] & ~x[1] & ~x[2] & ~x[11];
			partial_clause[2] 	= partial_clause_prev[2] & ~x[2];
			partial_clause[3] 	= partial_clause_prev[3] & ~x[11];
			partial_clause[4] 	= partial_clause_prev[4] & ~x[6] & ~x[7];
			partial_clause[5] 	= partial_clause_prev[5] & ~x[2];
			partial_clause[6] 	= partial_clause_prev[6] & ~x[2] & ~x[13];
			partial_clause[7] 	= partial_clause_prev[7] & ~x[2] & ~x[7];
			partial_clause[8] 	= partial_clause_prev[8] & ~x[2] & ~x[5] & ~x[11];
			partial_clause[9] 	= partial_clause_prev[9] & ~x[1] & ~x[2] & ~x[7] & ~x[8] & ~x[11] & ~x[12];
			partial_clause[10] 	= partial_clause_prev[10] & ~x[2] & ~x[10] & ~x[12];
			partial_clause[11] 	= partial_clause_prev[11] & ~x[2] & ~x[11] & ~x[12];
			partial_clause[12] 	= partial_clause_prev[12] & ~x[14];
			partial_clause[13] 	= partial_clause_prev[13] & ~x[3] & ~x[12];
			partial_clause[14] 	= partial_clause_prev[14] & 1'b1;
			partial_clause[15] 	= partial_clause_prev[15] & 1'b1;
			partial_clause[16] 	= partial_clause_prev[16] & ~x[4] & ~x[5] & ~x[13];
			partial_clause[17] 	= partial_clause_prev[17] & 1'b1;
			partial_clause[18] 	= partial_clause_prev[18] & 1'b1;
			partial_clause[19] 	= partial_clause_prev[19] & 1'b1;
			partial_clause[20] 	= partial_clause_prev[20] & ~x[15];
			partial_clause[21] 	= partial_clause_prev[21] & ~x[14];
			partial_clause[22] 	= partial_clause_prev[22] & ~x[8];
			partial_clause[23] 	= partial_clause_prev[23] & ~x[1] & ~x[2] & ~x[4] & ~x[6] & ~x[9] & ~x[11] & ~x[12] & ~x[13] & ~x[14];
			partial_clause[24] 	= partial_clause_prev[24] & ~x[1] & ~x[2] & ~x[3] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[11] & ~x[12] & ~x[15];
			partial_clause[25] 	= partial_clause_prev[25] & ~x[1] & ~x[9] & ~x[11] & ~x[12] & ~x[13];
			partial_clause[26] 	= partial_clause_prev[26] & 1'b1;
			partial_clause[27] 	= partial_clause_prev[27] & ~x[3] & ~x[9] & ~x[13];
			partial_clause[28] 	= partial_clause_prev[28] & ~x[1] & ~x[13];
			partial_clause[29] 	= partial_clause_prev[29] & ~x[7] & ~x[10] & ~x[15];
			partial_clause[30] 	= partial_clause_prev[30] & ~x[0] & ~x[15];
			partial_clause[31] 	= partial_clause_prev[31] & ~x[14];
			partial_clause[32] 	= partial_clause_prev[32] & 1'b1;
			partial_clause[33] 	= partial_clause_prev[33] & 1'b1;
			partial_clause[34] 	= partial_clause_prev[34] & 1'b1;
			partial_clause[35] 	= partial_clause_prev[35] & ~x[4] & ~x[8] & ~x[10] & ~x[11] & ~x[15];
			partial_clause[36] 	= partial_clause_prev[36] & ~x[5] & ~x[10];
			partial_clause[37] 	= partial_clause_prev[37] & ~x[8] & ~x[9];
			partial_clause[38] 	= partial_clause_prev[38] & ~x[5] & ~x[7];
			partial_clause[39] 	= partial_clause_prev[39] & 1'b1;
			partial_clause[40] 	= partial_clause_prev[40] & 1'b1;
			partial_clause[41] 	= partial_clause_prev[41] & 1'b1;
			partial_clause[42] 	= partial_clause_prev[42] & ~x[2];
			partial_clause[43] 	= partial_clause_prev[43] & ~x[10];
			partial_clause[44] 	= partial_clause_prev[44] & ~x[0] & ~x[10];
			partial_clause[45] 	= partial_clause_prev[45] & 1'b1;
			partial_clause[46] 	= partial_clause_prev[46] & ~x[0] & ~x[7] & ~x[9] & ~x[15];
			partial_clause[47] 	= partial_clause_prev[47] & 1'b1;
			partial_clause[48] 	= partial_clause_prev[48] & 1'b1;
			partial_clause[49] 	= partial_clause_prev[49] & 1'b1;
			partial_clause[50] 	= partial_clause_prev[50] & 1'b1;
			partial_clause[51] 	= partial_clause_prev[51] & 1'b1;
			partial_clause[52] 	= partial_clause_prev[52] & 1'b1;
			partial_clause[53] 	= partial_clause_prev[53] & 1'b1;
			partial_clause[54] 	= partial_clause_prev[54] & 1'b1;
			partial_clause[55] 	= partial_clause_prev[55] & 1'b1;
			partial_clause[56] 	= partial_clause_prev[56] & 1'b1;
			partial_clause[57] 	= partial_clause_prev[57] & ~x[0] & ~x[5];
			partial_clause[58] 	= partial_clause_prev[58] & ~x[9] & ~x[10];
			partial_clause[59] 	= partial_clause_prev[59] & ~x[6] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[14];
			partial_clause[60] 	= partial_clause_prev[60] & 1'b1;
			partial_clause[61] 	= partial_clause_prev[61] & ~x[8];
			partial_clause[62] 	= partial_clause_prev[62] & ~x[0] & ~x[1] & ~x[3] & ~x[7];
			partial_clause[63] 	= partial_clause_prev[63] & 1'b1;
			partial_clause[64] 	= partial_clause_prev[64] & 1'b1;
			partial_clause[65] 	= partial_clause_prev[65] & 1'b1;
			partial_clause[66] 	= partial_clause_prev[66] & 1'b1;
			partial_clause[67] 	= partial_clause_prev[67] & 1'b1;
			partial_clause[68] 	= partial_clause_prev[68] & ~x[0] & ~x[8] & ~x[10];
			partial_clause[69] 	= partial_clause_prev[69] & ~x[0] & ~x[7];
			partial_clause[70] 	= partial_clause_prev[70] & ~x[11];
			partial_clause[71] 	= partial_clause_prev[71] & ~x[5];
			partial_clause[72] 	= partial_clause_prev[72] & 1'b1;
			partial_clause[73] 	= partial_clause_prev[73] & ~x[5];
			partial_clause[74] 	= partial_clause_prev[74] & ~x[2] & ~x[12];
			partial_clause[75] 	= partial_clause_prev[75] & 1'b1;
			partial_clause[76] 	= partial_clause_prev[76] & ~x[5] & ~x[6] & ~x[13];
			partial_clause[77] 	= partial_clause_prev[77] & ~x[3] & ~x[15];
			partial_clause[78] 	= partial_clause_prev[78] & ~x[14];
			partial_clause[79] 	= partial_clause_prev[79] & 1'b1;
			partial_clause[80] 	= partial_clause_prev[80] & 1'b1;
			partial_clause[81] 	= partial_clause_prev[81] & 1'b1;
			partial_clause[82] 	= partial_clause_prev[82] & 1'b1;
			partial_clause[83] 	= partial_clause_prev[83] & 1'b1;
			partial_clause[84] 	= partial_clause_prev[84] & ~x[8] & ~x[9];
			partial_clause[85] 	= partial_clause_prev[85] & ~x[0] & ~x[7];
			partial_clause[86] 	= partial_clause_prev[86] & 1'b1;
			partial_clause[87] 	= partial_clause_prev[87] & ~x[15];
			partial_clause[88] 	= partial_clause_prev[88] & ~x[2];
			partial_clause[89] 	= partial_clause_prev[89] & 1'b1;
			partial_clause[90] 	= partial_clause_prev[90] & 1'b1;
			partial_clause[91] 	= partial_clause_prev[91] & 1'b1;
			partial_clause[92] 	= partial_clause_prev[92] & 1'b1;
			partial_clause[93] 	= partial_clause_prev[93] & ~x[2] & ~x[3] & ~x[4] & ~x[6] & ~x[7] & ~x[8] & ~x[11] & ~x[12] & ~x[13];
			partial_clause[94] 	= partial_clause_prev[94] & 1'b1;
			partial_clause[95] 	= partial_clause_prev[95] & ~x[12];
			partial_clause[96] 	= partial_clause_prev[96] & 1'b1;
			partial_clause[97] 	= partial_clause_prev[97] & ~x[0] & ~x[2] & ~x[8] & ~x[11] & ~x[12];
			partial_clause[98] 	= partial_clause_prev[98] & ~x[8] & ~x[10];
			partial_clause[99] 	= partial_clause_prev[99] & ~x[2] & ~x[3] & ~x[4] & ~x[5] & ~x[7] & ~x[10] & ~x[14] & ~x[15];
			partial_clause[100] 	= partial_clause_prev[100] & ~x[2];
			partial_clause[101] 	= partial_clause_prev[101] & 1'b1;
			partial_clause[102] 	= partial_clause_prev[102] & 1'b1;
			partial_clause[103] 	= partial_clause_prev[103] & ~x[3] & ~x[4] & ~x[12];
			partial_clause[104] 	= partial_clause_prev[104] & ~x[2] & ~x[7] & ~x[15];
			partial_clause[105] 	= partial_clause_prev[105] & ~x[9] & ~x[12] & ~x[14] & ~x[15];
			partial_clause[106] 	= partial_clause_prev[106] & 1'b1;
			partial_clause[107] 	= partial_clause_prev[107] & ~x[1] & ~x[10] & ~x[12];
			partial_clause[108] 	= partial_clause_prev[108] & ~x[2] & ~x[6] & ~x[9] & ~x[11] & ~x[13] & ~x[15];
			partial_clause[109] 	= partial_clause_prev[109] & 1'b1;
			partial_clause[110] 	= partial_clause_prev[110] & 1'b1;
			partial_clause[111] 	= partial_clause_prev[111] & 1'b1;
			partial_clause[112] 	= partial_clause_prev[112] & ~x[8];
			partial_clause[113] 	= partial_clause_prev[113] & 1'b1;
			partial_clause[114] 	= partial_clause_prev[114] & 1'b1;
			partial_clause[115] 	= partial_clause_prev[115] & ~x[6] & ~x[7] & ~x[9] & ~x[10] & ~x[11] & ~x[12] & ~x[13];
			partial_clause[116] 	= partial_clause_prev[116] & ~x[3] & ~x[5] & ~x[11] & ~x[15];
			partial_clause[117] 	= partial_clause_prev[117] & ~x[10];
			partial_clause[118] 	= partial_clause_prev[118] & ~x[2] & ~x[9];
			partial_clause[119] 	= partial_clause_prev[119] & ~x[2];
			partial_clause[120] 	= partial_clause_prev[120] & ~x[0] & ~x[3] & ~x[4] & ~x[5] & ~x[9] & ~x[10] & ~x[11] & ~x[15];
			partial_clause[121] 	= partial_clause_prev[121] & ~x[1] & ~x[3] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[11];
			partial_clause[122] 	= partial_clause_prev[122] & 1'b1;
			partial_clause[123] 	= partial_clause_prev[123] & ~x[0] & ~x[3] & ~x[6] & ~x[10] & ~x[11] & ~x[15];
			partial_clause[124] 	= partial_clause_prev[124] & 1'b1;
			partial_clause[125] 	= partial_clause_prev[125] & ~x[3];
			partial_clause[126] 	= partial_clause_prev[126] & 1'b1;
			partial_clause[127] 	= partial_clause_prev[127] & ~x[0] & ~x[1] & ~x[4] & ~x[5] & ~x[6] & ~x[7] & ~x[9] & ~x[11] & ~x[13] & ~x[14] & ~x[15];
			partial_clause[128] 	= partial_clause_prev[128] & 1'b1;
			partial_clause[129] 	= partial_clause_prev[129] & ~x[1] & ~x[3] & ~x[5] & ~x[11] & ~x[12] & ~x[15];
			partial_clause[130] 	= partial_clause_prev[130] & ~x[0];
			partial_clause[131] 	= partial_clause_prev[131] & 1'b1;
			partial_clause[132] 	= partial_clause_prev[132] & ~x[6] & ~x[9];
			partial_clause[133] 	= partial_clause_prev[133] & ~x[14];
			partial_clause[134] 	= partial_clause_prev[134] & ~x[0] & ~x[2] & ~x[3] & ~x[7] & ~x[9] & ~x[11] & ~x[12] & ~x[15];
			partial_clause[135] 	= partial_clause_prev[135] & ~x[9];
			partial_clause[136] 	= partial_clause_prev[136] & ~x[0] & ~x[2] & ~x[9] & ~x[11];
			partial_clause[137] 	= partial_clause_prev[137] & 1'b1;
			partial_clause[138] 	= partial_clause_prev[138] & 1'b1;
			partial_clause[139] 	= partial_clause_prev[139] & ~x[0] & ~x[5] & ~x[8] & ~x[9];
			partial_clause[140] 	= partial_clause_prev[140] & ~x[4] & ~x[7] & ~x[8] & ~x[11] & ~x[15];
			partial_clause[141] 	= partial_clause_prev[141] & 1'b1;
			partial_clause[142] 	= partial_clause_prev[142] & ~x[8] & ~x[10] & ~x[15];
			partial_clause[143] 	= partial_clause_prev[143] & 1'b1;
			partial_clause[144] 	= partial_clause_prev[144] & ~x[4] & ~x[6] & ~x[10] & ~x[12];
			partial_clause[145] 	= partial_clause_prev[145] & ~x[2];
			partial_clause[146] 	= partial_clause_prev[146] & ~x[1] & ~x[2] & ~x[8];
			partial_clause[147] 	= partial_clause_prev[147] & ~x[13];
			partial_clause[148] 	= partial_clause_prev[148] & ~x[7] & ~x[12];
			partial_clause[149] 	= partial_clause_prev[149] & 1'b1;
			partial_clause[150] 	= partial_clause_prev[150] & ~x[12];
			partial_clause[151] 	= partial_clause_prev[151] & 1'b1;
			partial_clause[152] 	= partial_clause_prev[152] & ~x[13];
			partial_clause[153] 	= partial_clause_prev[153] & ~x[2] & ~x[4];
			partial_clause[154] 	= partial_clause_prev[154] & ~x[9];
			partial_clause[155] 	= partial_clause_prev[155] & 1'b1;
			partial_clause[156] 	= partial_clause_prev[156] & ~x[7];
			partial_clause[157] 	= partial_clause_prev[157] & 1'b1;
			partial_clause[158] 	= partial_clause_prev[158] & ~x[0] & ~x[1] & ~x[2] & ~x[5] & ~x[7] & ~x[8] & ~x[9] & ~x[11] & ~x[12] & ~x[14];
			partial_clause[159] 	= partial_clause_prev[159] & ~x[3] & ~x[9];
			partial_clause[160] 	= partial_clause_prev[160] & 1'b1;
			partial_clause[161] 	= partial_clause_prev[161] & ~x[1] & ~x[6] & ~x[8] & ~x[12];
			partial_clause[162] 	= partial_clause_prev[162] & ~x[11];
			partial_clause[163] 	= partial_clause_prev[163] & 1'b1;
			partial_clause[164] 	= partial_clause_prev[164] & ~x[5] & ~x[8];
			partial_clause[165] 	= partial_clause_prev[165] & ~x[4] & ~x[9] & ~x[11];
			partial_clause[166] 	= partial_clause_prev[166] & ~x[8] & ~x[13];
			partial_clause[167] 	= partial_clause_prev[167] & 1'b1;
			partial_clause[168] 	= partial_clause_prev[168] & ~x[7];
			partial_clause[169] 	= partial_clause_prev[169] & 1'b1;
			partial_clause[170] 	= partial_clause_prev[170] & 1'b1;
			partial_clause[171] 	= partial_clause_prev[171] & ~x[2] & ~x[10] & ~x[11] & ~x[13];
			partial_clause[172] 	= partial_clause_prev[172] & 1'b1;
			partial_clause[173] 	= partial_clause_prev[173] & ~x[10];
			partial_clause[174] 	= partial_clause_prev[174] & ~x[5];
			partial_clause[175] 	= partial_clause_prev[175] & 1'b1;
			partial_clause[176] 	= partial_clause_prev[176] & 1'b1;
			partial_clause[177] 	= partial_clause_prev[177] & ~x[5] & ~x[13];
			partial_clause[178] 	= partial_clause_prev[178] & ~x[15];
			partial_clause[179] 	= partial_clause_prev[179] & 1'b1;
			partial_clause[180] 	= partial_clause_prev[180] & 1'b1;
			partial_clause[181] 	= partial_clause_prev[181] & 1'b1;
			partial_clause[182] 	= partial_clause_prev[182] & ~x[13];
			partial_clause[183] 	= partial_clause_prev[183] & ~x[5] & ~x[12] & ~x[13];
			partial_clause[184] 	= partial_clause_prev[184] & ~x[0] & ~x[1] & ~x[6] & ~x[8] & ~x[10];
			partial_clause[185] 	= partial_clause_prev[185] & ~x[1] & ~x[6] & ~x[14];
			partial_clause[186] 	= partial_clause_prev[186] & ~x[3] & ~x[5] & ~x[6];
			partial_clause[187] 	= partial_clause_prev[187] & 1'b1;
			partial_clause[188] 	= partial_clause_prev[188] & ~x[13];
			partial_clause[189] 	= partial_clause_prev[189] & 1'b1;
			partial_clause[190] 	= partial_clause_prev[190] & ~x[14];
			partial_clause[191] 	= partial_clause_prev[191] & ~x[7];
			partial_clause[192] 	= partial_clause_prev[192] & ~x[15];
			partial_clause[193] 	= partial_clause_prev[193] & 1'b1;
			partial_clause[194] 	= partial_clause_prev[194] & ~x[9];
			partial_clause[195] 	= partial_clause_prev[195] & ~x[4] & ~x[7] & ~x[14] & ~x[15];
			partial_clause[196] 	= partial_clause_prev[196] & ~x[1];
			partial_clause[197] 	= partial_clause_prev[197] & ~x[6];
			partial_clause[198] 	= partial_clause_prev[198] & 1'b1;
			partial_clause[199] 	= partial_clause_prev[199] & 1'b1;
			partial_clause[200] 	= partial_clause_prev[200] & ~x[6];
			partial_clause[201] 	= partial_clause_prev[201] & ~x[2] & ~x[4] & ~x[6] & ~x[12];
			partial_clause[202] 	= partial_clause_prev[202] & ~x[12] & ~x[13];
			partial_clause[203] 	= partial_clause_prev[203] & ~x[2];
			partial_clause[204] 	= partial_clause_prev[204] & ~x[1] & ~x[3] & ~x[4] & ~x[5] & ~x[7] & ~x[11];
			partial_clause[205] 	= partial_clause_prev[205] & 1'b1;
			partial_clause[206] 	= partial_clause_prev[206] & ~x[6] & ~x[8];
			partial_clause[207] 	= partial_clause_prev[207] & ~x[15];
			partial_clause[208] 	= partial_clause_prev[208] & ~x[2] & ~x[13];
			partial_clause[209] 	= partial_clause_prev[209] & 1'b1;
			partial_clause[210] 	= partial_clause_prev[210] & ~x[1] & ~x[3];
			partial_clause[211] 	= partial_clause_prev[211] & 1'b1;
			partial_clause[212] 	= partial_clause_prev[212] & 1'b1;
			partial_clause[213] 	= partial_clause_prev[213] & 1'b1;
			partial_clause[214] 	= partial_clause_prev[214] & 1'b1;
			partial_clause[215] 	= partial_clause_prev[215] & 1'b1;
			partial_clause[216] 	= partial_clause_prev[216] & 1'b1;
			partial_clause[217] 	= partial_clause_prev[217] & ~x[3] & ~x[5];
			partial_clause[218] 	= partial_clause_prev[218] & ~x[9];
			partial_clause[219] 	= partial_clause_prev[219] & 1'b1;
			partial_clause[220] 	= partial_clause_prev[220] & ~x[0] & ~x[10];
			partial_clause[221] 	= partial_clause_prev[221] & 1'b1;
			partial_clause[222] 	= partial_clause_prev[222] & 1'b1;
			partial_clause[223] 	= partial_clause_prev[223] & 1'b1;
			partial_clause[224] 	= partial_clause_prev[224] & ~x[0] & ~x[1] & ~x[6];
			partial_clause[225] 	= partial_clause_prev[225] & ~x[4] & ~x[8] & ~x[13];
			partial_clause[226] 	= partial_clause_prev[226] & ~x[1] & ~x[2] & ~x[5] & ~x[13] & ~x[15];
			partial_clause[227] 	= partial_clause_prev[227] & 1'b1;
			partial_clause[228] 	= partial_clause_prev[228] & ~x[8] & ~x[15];
			partial_clause[229] 	= partial_clause_prev[229] & ~x[1];
			partial_clause[230] 	= partial_clause_prev[230] & ~x[0] & ~x[1] & ~x[2] & ~x[3] & ~x[8] & ~x[9] & ~x[13];
			partial_clause[231] 	= partial_clause_prev[231] & 1'b1;
			partial_clause[232] 	= partial_clause_prev[232] & 1'b1;
			partial_clause[233] 	= partial_clause_prev[233] & ~x[5];
			partial_clause[234] 	= partial_clause_prev[234] & ~x[14];
			partial_clause[235] 	= partial_clause_prev[235] & 1'b1;
			partial_clause[236] 	= partial_clause_prev[236] & 1'b1;
			partial_clause[237] 	= partial_clause_prev[237] & ~x[2];
			partial_clause[238] 	= partial_clause_prev[238] & ~x[6];
			partial_clause[239] 	= partial_clause_prev[239] & 1'b1;
			partial_clause[240] 	= partial_clause_prev[240] & ~x[13];
			partial_clause[241] 	= partial_clause_prev[241] & 1'b1;
			partial_clause[242] 	= partial_clause_prev[242] & ~x[6] & ~x[10];
			partial_clause[243] 	= partial_clause_prev[243] & ~x[2] & ~x[4] & ~x[8] & ~x[10];
			partial_clause[244] 	= partial_clause_prev[244] & ~x[15];
			partial_clause[245] 	= partial_clause_prev[245] & 1'b1;
			partial_clause[246] 	= partial_clause_prev[246] & 1'b1;
			partial_clause[247] 	= partial_clause_prev[247] & ~x[0] & ~x[1] & ~x[4] & ~x[11] & ~x[13] & ~x[14];
			partial_clause[248] 	= partial_clause_prev[248] & ~x[0] & ~x[3] & ~x[4] & ~x[5] & ~x[6] & ~x[10] & ~x[12] & ~x[14] & ~x[15];
			partial_clause[249] 	= partial_clause_prev[249] & ~x[13] & ~x[14];
			partial_clause[250] 	= partial_clause_prev[250] & ~x[4] & ~x[5] & ~x[6] & ~x[9] & ~x[11] & ~x[12] & ~x[14];
			partial_clause[251] 	= partial_clause_prev[251] & 1'b1;
			partial_clause[252] 	= partial_clause_prev[252] & ~x[1] & ~x[5] & ~x[7] & ~x[13] & ~x[14];
			partial_clause[253] 	= partial_clause_prev[253] & ~x[5];
			partial_clause[254] 	= partial_clause_prev[254] & ~x[4];
			partial_clause[255] 	= partial_clause_prev[255] & ~x[13];
			partial_clause[256] 	= partial_clause_prev[256] & 1'b1;
			partial_clause[257] 	= partial_clause_prev[257] & ~x[3] & ~x[5];
			partial_clause[258] 	= partial_clause_prev[258] & ~x[1] & ~x[6] & ~x[8];
			partial_clause[259] 	= partial_clause_prev[259] & 1'b1;
			partial_clause[260] 	= partial_clause_prev[260] & ~x[2] & ~x[3];
			partial_clause[261] 	= partial_clause_prev[261] & ~x[6] & ~x[12];
			partial_clause[262] 	= partial_clause_prev[262] & ~x[6] & ~x[9] & ~x[11];
			partial_clause[263] 	= partial_clause_prev[263] & ~x[1];
			partial_clause[264] 	= partial_clause_prev[264] & ~x[9];
			partial_clause[265] 	= partial_clause_prev[265] & 1'b1;
			partial_clause[266] 	= partial_clause_prev[266] & ~x[6] & ~x[8];
			partial_clause[267] 	= partial_clause_prev[267] & ~x[6] & ~x[8];
			partial_clause[268] 	= partial_clause_prev[268] & ~x[1] & ~x[2] & ~x[4] & ~x[8] & ~x[10];
			partial_clause[269] 	= partial_clause_prev[269] & ~x[0] & ~x[1] & ~x[5] & ~x[8] & ~x[9] & ~x[11] & ~x[13];
			partial_clause[270] 	= partial_clause_prev[270] & 1'b1;
			partial_clause[271] 	= partial_clause_prev[271] & 1'b1;
			partial_clause[272] 	= partial_clause_prev[272] & ~x[4] & ~x[13];
			partial_clause[273] 	= partial_clause_prev[273] & ~x[0] & ~x[1] & ~x[6] & ~x[8] & ~x[9] & ~x[10] & ~x[11];
			partial_clause[274] 	= partial_clause_prev[274] & ~x[1] & ~x[12];
			partial_clause[275] 	= partial_clause_prev[275] & 1'b1;
			partial_clause[276] 	= partial_clause_prev[276] & ~x[15];
			partial_clause[277] 	= partial_clause_prev[277] & ~x[15];
			partial_clause[278] 	= partial_clause_prev[278] & 1'b1;
			partial_clause[279] 	= partial_clause_prev[279] & ~x[1] & ~x[4] & ~x[11] & ~x[13] & ~x[14];
			partial_clause[280] 	= partial_clause_prev[280] & 1'b1;
			partial_clause[281] 	= partial_clause_prev[281] & ~x[0] & ~x[13];
			partial_clause[282] 	= partial_clause_prev[282] & ~x[14];
			partial_clause[283] 	= partial_clause_prev[283] & ~x[7];
			partial_clause[284] 	= partial_clause_prev[284] & 1'b1;
			partial_clause[285] 	= partial_clause_prev[285] & 1'b1;
			partial_clause[286] 	= partial_clause_prev[286] & 1'b1;
			partial_clause[287] 	= partial_clause_prev[287] & ~x[0] & ~x[1] & ~x[6] & ~x[8] & ~x[12] & ~x[13] & ~x[14] & ~x[15];
			partial_clause[288] 	= partial_clause_prev[288] & 1'b1;
			partial_clause[289] 	= partial_clause_prev[289] & ~x[2] & ~x[3];
			partial_clause[290] 	= partial_clause_prev[290] & ~x[9] & ~x[14];
			partial_clause[291] 	= partial_clause_prev[291] & 1'b1;
			partial_clause[292] 	= partial_clause_prev[292] & ~x[5] & ~x[12];
			partial_clause[293] 	= partial_clause_prev[293] & ~x[0];
			partial_clause[294] 	= partial_clause_prev[294] & 1'b1;
			partial_clause[295] 	= partial_clause_prev[295] & 1'b1;
			partial_clause[296] 	= partial_clause_prev[296] & 1'b1;
			partial_clause[297] 	= partial_clause_prev[297] & ~x[2];
			partial_clause[298] 	= partial_clause_prev[298] & 1'b1;
			partial_clause[299] 	= partial_clause_prev[299] & 1'b1;
			partial_clause[300] 	= partial_clause_prev[300] & 1'b1;
			partial_clause[301] 	= partial_clause_prev[301] & ~x[2] & ~x[5] & ~x[6];
			partial_clause[302] 	= partial_clause_prev[302] & ~x[4];
			partial_clause[303] 	= partial_clause_prev[303] & 1'b1;
			partial_clause[304] 	= partial_clause_prev[304] & ~x[8];
			partial_clause[305] 	= partial_clause_prev[305] & ~x[7];
			partial_clause[306] 	= partial_clause_prev[306] & ~x[13];
			partial_clause[307] 	= partial_clause_prev[307] & ~x[6];
			partial_clause[308] 	= partial_clause_prev[308] & ~x[3] & ~x[9] & ~x[11] & ~x[13];
			partial_clause[309] 	= partial_clause_prev[309] & ~x[7] & ~x[10];
			partial_clause[310] 	= partial_clause_prev[310] & 1'b1;
			partial_clause[311] 	= partial_clause_prev[311] & ~x[5] & ~x[7];
			partial_clause[312] 	= partial_clause_prev[312] & 1'b1;
			partial_clause[313] 	= partial_clause_prev[313] & ~x[6];
			partial_clause[314] 	= partial_clause_prev[314] & 1'b1;
			partial_clause[315] 	= partial_clause_prev[315] & 1'b1;
			partial_clause[316] 	= partial_clause_prev[316] & ~x[0] & ~x[1] & ~x[5] & ~x[7] & ~x[10];
			partial_clause[317] 	= partial_clause_prev[317] & ~x[4] & ~x[6] & ~x[13] & ~x[15];
			partial_clause[318] 	= partial_clause_prev[318] & 1'b1;
			partial_clause[319] 	= partial_clause_prev[319] & 1'b1;
			partial_clause[320] 	= partial_clause_prev[320] & ~x[2];
			partial_clause[321] 	= partial_clause_prev[321] & ~x[9];
			partial_clause[322] 	= partial_clause_prev[322] & ~x[2];
			partial_clause[323] 	= partial_clause_prev[323] & ~x[12];
			partial_clause[324] 	= partial_clause_prev[324] & 1'b1;
			partial_clause[325] 	= partial_clause_prev[325] & ~x[0] & ~x[1] & ~x[3] & ~x[5] & ~x[6] & ~x[7] & ~x[8] & ~x[9] & ~x[12] & ~x[13] & ~x[14];
			partial_clause[326] 	= partial_clause_prev[326] & ~x[10] & ~x[13];
			partial_clause[327] 	= partial_clause_prev[327] & ~x[0];
			partial_clause[328] 	= partial_clause_prev[328] & ~x[1];
			partial_clause[329] 	= partial_clause_prev[329] & 1'b1;
			partial_clause[330] 	= partial_clause_prev[330] & ~x[4] & ~x[10] & ~x[15];
			partial_clause[331] 	= partial_clause_prev[331] & 1'b1;
			partial_clause[332] 	= partial_clause_prev[332] & ~x[14];
			partial_clause[333] 	= partial_clause_prev[333] & ~x[8];
			partial_clause[334] 	= partial_clause_prev[334] & ~x[0] & ~x[1] & ~x[15];
			partial_clause[335] 	= partial_clause_prev[335] & 1'b1;
			partial_clause[336] 	= partial_clause_prev[336] & 1'b1;
			partial_clause[337] 	= partial_clause_prev[337] & ~x[12] & ~x[13] & ~x[15];
			partial_clause[338] 	= partial_clause_prev[338] & 1'b1;
			partial_clause[339] 	= partial_clause_prev[339] & ~x[2] & ~x[4] & ~x[10];
			partial_clause[340] 	= partial_clause_prev[340] & ~x[5] & ~x[12] & ~x[15];
			partial_clause[341] 	= partial_clause_prev[341] & 1'b1;
			partial_clause[342] 	= partial_clause_prev[342] & ~x[2] & ~x[3] & ~x[15];
			partial_clause[343] 	= partial_clause_prev[343] & ~x[0] & ~x[7] & ~x[9] & ~x[12] & ~x[14];
			partial_clause[344] 	= partial_clause_prev[344] & ~x[2] & ~x[10];
			partial_clause[345] 	= partial_clause_prev[345] & 1'b1;
			partial_clause[346] 	= partial_clause_prev[346] & ~x[3] & ~x[4] & ~x[9];
			partial_clause[347] 	= partial_clause_prev[347] & ~x[4] & ~x[5] & ~x[9];
			partial_clause[348] 	= partial_clause_prev[348] & ~x[2];
			partial_clause[349] 	= partial_clause_prev[349] & 1'b1;
			partial_clause[350] 	= partial_clause_prev[350] & ~x[5] & ~x[7] & ~x[8] & ~x[10] & ~x[12] & ~x[14];
			partial_clause[351] 	= partial_clause_prev[351] & 1'b1;
			partial_clause[352] 	= partial_clause_prev[352] & 1'b1;
			partial_clause[353] 	= partial_clause_prev[353] & 1'b1;
			partial_clause[354] 	= partial_clause_prev[354] & ~x[3] & ~x[11];
			partial_clause[355] 	= partial_clause_prev[355] & 1'b1;
			partial_clause[356] 	= partial_clause_prev[356] & 1'b1;
			partial_clause[357] 	= partial_clause_prev[357] & 1'b1;
			partial_clause[358] 	= partial_clause_prev[358] & ~x[0] & ~x[2];
			partial_clause[359] 	= partial_clause_prev[359] & ~x[7];
			partial_clause[360] 	= partial_clause_prev[360] & ~x[1] & ~x[2] & ~x[10] & ~x[11] & ~x[12] & ~x[15];
			partial_clause[361] 	= partial_clause_prev[361] & ~x[1] & ~x[10];
			partial_clause[362] 	= partial_clause_prev[362] & ~x[3];
			partial_clause[363] 	= partial_clause_prev[363] & ~x[0] & ~x[1] & ~x[3] & ~x[11] & ~x[13] & ~x[14];
			partial_clause[364] 	= partial_clause_prev[364] & 1'b1;
			partial_clause[365] 	= partial_clause_prev[365] & ~x[2];
			partial_clause[366] 	= partial_clause_prev[366] & ~x[2] & ~x[7] & ~x[11];
			partial_clause[367] 	= partial_clause_prev[367] & ~x[12];
			partial_clause[368] 	= partial_clause_prev[368] & 1'b1;
			partial_clause[369] 	= partial_clause_prev[369] & ~x[4] & ~x[10];
			partial_clause[370] 	= partial_clause_prev[370] & ~x[0] & ~x[15];
			partial_clause[371] 	= partial_clause_prev[371] & 1'b1;
			partial_clause[372] 	= partial_clause_prev[372] & ~x[1] & ~x[2] & ~x[9];
			partial_clause[373] 	= partial_clause_prev[373] & 1'b1;
			partial_clause[374] 	= partial_clause_prev[374] & 1'b1;
			partial_clause[375] 	= partial_clause_prev[375] & 1'b1;
			partial_clause[376] 	= partial_clause_prev[376] & 1'b1;
			partial_clause[377] 	= partial_clause_prev[377] & ~x[8] & ~x[9] & ~x[11];
			partial_clause[378] 	= partial_clause_prev[378] & ~x[13];
			partial_clause[379] 	= partial_clause_prev[379] & ~x[0] & ~x[6] & ~x[15];
			partial_clause[380] 	= partial_clause_prev[380] & 1'b1;
			partial_clause[381] 	= partial_clause_prev[381] & ~x[0] & ~x[2] & ~x[10] & ~x[13];
			partial_clause[382] 	= partial_clause_prev[382] & 1'b1;
			partial_clause[383] 	= partial_clause_prev[383] & 1'b1;
			partial_clause[384] 	= partial_clause_prev[384] & 1'b1;
			partial_clause[385] 	= partial_clause_prev[385] & ~x[4];
			partial_clause[386] 	= partial_clause_prev[386] & 1'b1;
			partial_clause[387] 	= partial_clause_prev[387] & ~x[0] & ~x[2] & ~x[7] & ~x[12] & ~x[14];
			partial_clause[388] 	= partial_clause_prev[388] & ~x[1] & ~x[3] & ~x[14];
			partial_clause[389] 	= partial_clause_prev[389] & 1'b1;
			partial_clause[390] 	= partial_clause_prev[390] & ~x[0] & ~x[2] & ~x[3] & ~x[9];
			partial_clause[391] 	= partial_clause_prev[391] & 1'b1;
			partial_clause[392] 	= partial_clause_prev[392] & 1'b1;
			partial_clause[393] 	= partial_clause_prev[393] & 1'b1;
			partial_clause[394] 	= partial_clause_prev[394] & 1'b1;
			partial_clause[395] 	= partial_clause_prev[395] & ~x[9];
			partial_clause[396] 	= partial_clause_prev[396] & 1'b1;
			partial_clause[397] 	= partial_clause_prev[397] & 1'b1;
			partial_clause[398] 	= partial_clause_prev[398] & 1'b1;
			partial_clause[399] 	= partial_clause_prev[399] & ~x[3];
			partial_clause[400] 	= partial_clause_prev[400] & ~x[3] & ~x[4] & ~x[10];
			partial_clause[401] 	= partial_clause_prev[401] & ~x[3] & ~x[13] & ~x[15];
			partial_clause[402] 	= partial_clause_prev[402] & ~x[0] & ~x[12] & ~x[14];
			partial_clause[403] 	= partial_clause_prev[403] & ~x[5] & ~x[9];
			partial_clause[404] 	= partial_clause_prev[404] & 1'b1;
			partial_clause[405] 	= partial_clause_prev[405] & ~x[10];
			partial_clause[406] 	= partial_clause_prev[406] & ~x[7];
			partial_clause[407] 	= partial_clause_prev[407] & ~x[0] & ~x[9];
			partial_clause[408] 	= partial_clause_prev[408] & 1'b1;
			partial_clause[409] 	= partial_clause_prev[409] & ~x[1] & ~x[2] & ~x[5] & ~x[6] & ~x[7] & ~x[10] & ~x[11] & ~x[13] & ~x[14];
			partial_clause[410] 	= partial_clause_prev[410] & ~x[13];
			partial_clause[411] 	= partial_clause_prev[411] & 1'b1;
			partial_clause[412] 	= partial_clause_prev[412] & ~x[4] & ~x[14];
			partial_clause[413] 	= partial_clause_prev[413] & ~x[8] & ~x[15];
			partial_clause[414] 	= partial_clause_prev[414] & ~x[3] & ~x[12];
			partial_clause[415] 	= partial_clause_prev[415] & ~x[6];
			partial_clause[416] 	= partial_clause_prev[416] & ~x[3] & ~x[7] & ~x[14];
			partial_clause[417] 	= partial_clause_prev[417] & ~x[5] & ~x[8] & ~x[15];
			partial_clause[418] 	= partial_clause_prev[418] & ~x[6] & ~x[9] & ~x[12] & ~x[14];
			partial_clause[419] 	= partial_clause_prev[419] & 1'b1;
			partial_clause[420] 	= partial_clause_prev[420] & 1'b1;
			partial_clause[421] 	= partial_clause_prev[421] & ~x[2] & ~x[13] & ~x[15];
			partial_clause[422] 	= partial_clause_prev[422] & ~x[0] & ~x[11];
			partial_clause[423] 	= partial_clause_prev[423] & 1'b1;
			partial_clause[424] 	= partial_clause_prev[424] & 1'b1;
			partial_clause[425] 	= partial_clause_prev[425] & ~x[5] & ~x[9];
			partial_clause[426] 	= partial_clause_prev[426] & ~x[2] & ~x[8] & ~x[10] & ~x[14] & ~x[15];
			partial_clause[427] 	= partial_clause_prev[427] & ~x[6];
			partial_clause[428] 	= partial_clause_prev[428] & 1'b1;
			partial_clause[429] 	= partial_clause_prev[429] & 1'b1;
			partial_clause[430] 	= partial_clause_prev[430] & ~x[3] & ~x[14];
			partial_clause[431] 	= partial_clause_prev[431] & ~x[3];
			partial_clause[432] 	= partial_clause_prev[432] & ~x[0] & ~x[1] & ~x[3] & ~x[8] & ~x[9] & ~x[12] & ~x[14];
			partial_clause[433] 	= partial_clause_prev[433] & ~x[11];
			partial_clause[434] 	= partial_clause_prev[434] & 1'b1;
			partial_clause[435] 	= partial_clause_prev[435] & ~x[1] & ~x[3] & ~x[8] & ~x[9] & ~x[11] & ~x[12];
			partial_clause[436] 	= partial_clause_prev[436] & ~x[11];
			partial_clause[437] 	= partial_clause_prev[437] & ~x[5] & ~x[8] & ~x[9];
			partial_clause[438] 	= partial_clause_prev[438] & 1'b1;
			partial_clause[439] 	= partial_clause_prev[439] & ~x[0] & ~x[2] & ~x[5] & ~x[10];
			partial_clause[440] 	= partial_clause_prev[440] & 1'b1;
			partial_clause[441] 	= partial_clause_prev[441] & ~x[3];
			partial_clause[442] 	= partial_clause_prev[442] & 1'b1;
			partial_clause[443] 	= partial_clause_prev[443] & ~x[8] & ~x[11] & ~x[12];
			partial_clause[444] 	= partial_clause_prev[444] & 1'b1;
			partial_clause[445] 	= partial_clause_prev[445] & 1'b1;
			partial_clause[446] 	= partial_clause_prev[446] & ~x[2] & ~x[4] & ~x[13];
			partial_clause[447] 	= partial_clause_prev[447] & ~x[1] & ~x[9] & ~x[14];
			partial_clause[448] 	= partial_clause_prev[448] & 1'b1;
			partial_clause[449] 	= partial_clause_prev[449] & ~x[2];
			partial_clause[450] 	= partial_clause_prev[450] & ~x[15];
			partial_clause[451] 	= partial_clause_prev[451] & 1'b1;
			partial_clause[452] 	= partial_clause_prev[452] & ~x[2] & ~x[13];
			partial_clause[453] 	= partial_clause_prev[453] & ~x[10];
			partial_clause[454] 	= partial_clause_prev[454] & 1'b1;
			partial_clause[455] 	= partial_clause_prev[455] & ~x[4] & ~x[9] & ~x[10];
			partial_clause[456] 	= partial_clause_prev[456] & ~x[2] & ~x[4] & ~x[9] & ~x[14];
			partial_clause[457] 	= partial_clause_prev[457] & 1'b1;
			partial_clause[458] 	= partial_clause_prev[458] & ~x[1] & ~x[3] & ~x[15];
			partial_clause[459] 	= partial_clause_prev[459] & ~x[9];
			partial_clause[460] 	= partial_clause_prev[460] & ~x[5] & ~x[9];
			partial_clause[461] 	= partial_clause_prev[461] & ~x[1];
			partial_clause[462] 	= partial_clause_prev[462] & ~x[14];
			partial_clause[463] 	= partial_clause_prev[463] & 1'b1;
			partial_clause[464] 	= partial_clause_prev[464] & ~x[5];
			partial_clause[465] 	= partial_clause_prev[465] & ~x[8] & ~x[13];
			partial_clause[466] 	= partial_clause_prev[466] & ~x[6] & ~x[7] & ~x[10];
			partial_clause[467] 	= partial_clause_prev[467] & ~x[3];
			partial_clause[468] 	= partial_clause_prev[468] & ~x[0] & ~x[1];
			partial_clause[469] 	= partial_clause_prev[469] & ~x[1] & ~x[3] & ~x[4] & ~x[11] & ~x[12] & ~x[15];
			partial_clause[470] 	= partial_clause_prev[470] & 1'b1;
			partial_clause[471] 	= partial_clause_prev[471] & ~x[2] & ~x[5];
			partial_clause[472] 	= partial_clause_prev[472] & ~x[10];
			partial_clause[473] 	= partial_clause_prev[473] & ~x[5] & ~x[14];
			partial_clause[474] 	= partial_clause_prev[474] & 1'b1;
			partial_clause[475] 	= partial_clause_prev[475] & ~x[9] & ~x[10];
			partial_clause[476] 	= partial_clause_prev[476] & ~x[12];
			partial_clause[477] 	= partial_clause_prev[477] & ~x[9] & ~x[13];
			partial_clause[478] 	= partial_clause_prev[478] & ~x[3] & ~x[7] & ~x[8] & ~x[13];
			partial_clause[479] 	= partial_clause_prev[479] & 1'b1;
			partial_clause[480] 	= partial_clause_prev[480] & ~x[1] & ~x[2] & ~x[3] & ~x[6] & ~x[10] & ~x[11] & ~x[12] & ~x[13] & ~x[15];
			partial_clause[481] 	= partial_clause_prev[481] & 1'b1;
			partial_clause[482] 	= partial_clause_prev[482] & ~x[1] & ~x[14];
			partial_clause[483] 	= partial_clause_prev[483] & ~x[0];
			partial_clause[484] 	= partial_clause_prev[484] & ~x[5];
			partial_clause[485] 	= partial_clause_prev[485] & 1'b1;
			partial_clause[486] 	= partial_clause_prev[486] & ~x[1] & ~x[3] & ~x[8] & ~x[11] & ~x[13];
			partial_clause[487] 	= partial_clause_prev[487] & ~x[10] & ~x[14];
			partial_clause[488] 	= partial_clause_prev[488] & 1'b1;
			partial_clause[489] 	= partial_clause_prev[489] & 1'b1;
			partial_clause[490] 	= partial_clause_prev[490] & 1'b1;
			partial_clause[491] 	= partial_clause_prev[491] & 1'b1;
			partial_clause[492] 	= partial_clause_prev[492] & ~x[2] & ~x[3] & ~x[13];
			partial_clause[493] 	= partial_clause_prev[493] & 1'b1;
			partial_clause[494] 	= partial_clause_prev[494] & 1'b1;
			partial_clause[495] 	= partial_clause_prev[495] & ~x[9] & ~x[12];
			partial_clause[496] 	= partial_clause_prev[496] & 1'b1;
			partial_clause[497] 	= partial_clause_prev[497] & 1'b1;
			partial_clause[498] 	= partial_clause_prev[498] & 1'b1;
			partial_clause[499] 	= partial_clause_prev[499] & 1'b1;
		end
	end
endmodule


